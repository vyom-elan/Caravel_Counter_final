magic
tech sky130A
magscale 1 2
timestamp 1706777037
<< checkpaint >>
rect -12658 -11586 596582 715522
<< metal1 >>
rect 35986 2864 35992 2916
rect 36044 2904 36050 2916
rect 40402 2904 40408 2916
rect 36044 2876 40408 2904
rect 36044 2864 36050 2876
rect 40402 2864 40408 2876
rect 40460 2864 40466 2916
rect 134334 2864 134340 2916
rect 134392 2904 134398 2916
rect 145144 2904 145150 2916
rect 134392 2876 145150 2904
rect 134392 2864 134398 2876
rect 145144 2864 145150 2876
rect 145202 2864 145208 2916
rect 169570 2864 169576 2916
rect 169628 2904 169634 2916
rect 178264 2904 178270 2916
rect 169628 2876 178270 2904
rect 169628 2864 169634 2876
rect 178264 2864 178270 2876
rect 178322 2864 178328 2916
rect 359320 2864 359326 2916
rect 359378 2904 359384 2916
rect 363322 2904 363328 2916
rect 359378 2876 363328 2904
rect 359378 2864 359384 2876
rect 363322 2864 363328 2876
rect 363380 2864 363386 2916
rect 364058 2864 364064 2916
rect 364116 2904 364122 2916
rect 365714 2904 365720 2916
rect 364116 2876 365720 2904
rect 364116 2864 364122 2876
rect 365714 2864 365720 2876
rect 365772 2864 365778 2916
rect 365944 2864 365950 2916
rect 366002 2904 366008 2916
rect 370038 2904 370044 2916
rect 366002 2876 370044 2904
rect 366002 2864 366008 2876
rect 370038 2864 370044 2876
rect 370096 2864 370102 2916
rect 370360 2864 370366 2916
rect 370418 2904 370424 2916
rect 375190 2904 375196 2916
rect 370418 2876 375196 2904
rect 370418 2864 370424 2876
rect 375190 2864 375196 2876
rect 375248 2864 375254 2916
rect 376984 2864 376990 2916
rect 377042 2904 377048 2916
rect 382274 2904 382280 2916
rect 377042 2876 382280 2904
rect 377042 2864 377048 2876
rect 382274 2864 382280 2876
rect 382332 2864 382338 2916
rect 385816 2864 385822 2916
rect 385874 2904 385880 2916
rect 391842 2904 391848 2916
rect 385874 2876 391848 2904
rect 385874 2864 385880 2876
rect 391842 2864 391848 2876
rect 391900 2864 391906 2916
rect 393222 2864 393228 2916
rect 393280 2904 393286 2916
rect 394050 2904 394056 2916
rect 393280 2876 394056 2904
rect 393280 2864 393286 2876
rect 394050 2864 394056 2876
rect 394108 2864 394114 2916
rect 394648 2864 394654 2916
rect 394706 2904 394712 2916
rect 400858 2904 400864 2916
rect 394706 2876 400864 2904
rect 394706 2864 394712 2876
rect 400858 2864 400864 2876
rect 400916 2864 400922 2916
rect 30098 2796 30104 2848
rect 30156 2836 30162 2848
rect 37182 2836 37188 2848
rect 30156 2808 37188 2836
rect 30156 2796 30162 2808
rect 37182 2796 37188 2808
rect 37240 2796 37246 2848
rect 41874 2796 41880 2848
rect 41932 2836 41938 2848
rect 49602 2836 49608 2848
rect 41932 2808 49608 2836
rect 41932 2796 41938 2808
rect 49602 2796 49608 2808
rect 49660 2796 49666 2848
rect 51350 2796 51356 2848
rect 51408 2836 51414 2848
rect 59262 2836 59268 2848
rect 51408 2808 59268 2836
rect 51408 2796 51414 2808
rect 59262 2796 59268 2808
rect 59320 2796 59326 2848
rect 60826 2796 60832 2848
rect 60884 2836 60890 2848
rect 68922 2836 68928 2848
rect 60884 2808 68928 2836
rect 60884 2796 60890 2808
rect 68922 2796 68928 2808
rect 68980 2796 68986 2848
rect 70302 2796 70308 2848
rect 70360 2836 70366 2848
rect 77202 2836 77208 2848
rect 70360 2808 77208 2836
rect 70360 2796 70366 2808
rect 77202 2796 77208 2808
rect 77260 2796 77266 2848
rect 82078 2796 82084 2848
rect 82136 2836 82142 2848
rect 96568 2836 96574 2848
rect 82136 2808 96574 2836
rect 82136 2796 82142 2808
rect 96568 2796 96574 2808
rect 96626 2796 96632 2848
rect 153010 2796 153016 2848
rect 153068 2836 153074 2848
rect 162808 2836 162814 2848
rect 153068 2808 162814 2836
rect 153068 2796 153074 2808
rect 162808 2796 162814 2808
rect 162866 2796 162872 2848
rect 351592 2796 351598 2848
rect 351650 2836 351656 2848
rect 355042 2836 355048 2848
rect 351650 2808 355048 2836
rect 351650 2796 351656 2808
rect 355042 2796 355048 2808
rect 355100 2796 355106 2848
rect 358216 2796 358222 2848
rect 358274 2836 358280 2848
rect 361666 2836 361672 2848
rect 358274 2808 361672 2836
rect 358274 2796 358280 2808
rect 361666 2796 361672 2808
rect 361724 2796 361730 2848
rect 367048 2796 367054 2848
rect 367106 2836 367112 2848
rect 371234 2836 371240 2848
rect 367106 2808 371240 2836
rect 367106 2796 367112 2808
rect 371234 2796 371240 2808
rect 371292 2796 371298 2848
rect 371326 2796 371332 2848
rect 371384 2836 371390 2848
rect 373994 2836 374000 2848
rect 371384 2808 374000 2836
rect 371384 2796 371390 2808
rect 373994 2796 374000 2808
rect 374052 2796 374058 2848
rect 375880 2796 375886 2848
rect 375938 2836 375944 2848
rect 380894 2836 380900 2848
rect 375938 2808 380900 2836
rect 375938 2796 375944 2808
rect 380894 2796 380900 2808
rect 380952 2796 380958 2848
rect 389128 2796 389134 2848
rect 389186 2836 389192 2848
rect 393498 2836 393504 2848
rect 389186 2808 393504 2836
rect 389186 2796 389192 2808
rect 393498 2796 393504 2808
rect 393556 2796 393562 2848
rect 395752 2796 395758 2848
rect 395810 2836 395816 2848
rect 402330 2836 402336 2848
rect 395810 2808 402336 2836
rect 395810 2796 395816 2808
rect 402330 2796 402336 2808
rect 402388 2796 402394 2848
rect 404584 2796 404590 2848
rect 404642 2836 404648 2848
rect 411714 2836 411720 2848
rect 404642 2808 411720 2836
rect 404642 2796 404648 2808
rect 411714 2796 411720 2808
rect 411772 2796 411778 2848
rect 449848 2796 449854 2848
rect 449906 2836 449912 2848
rect 460382 2836 460388 2848
rect 449906 2808 460388 2836
rect 449906 2796 449912 2808
rect 460382 2796 460388 2808
rect 460440 2796 460446 2848
rect 478874 2796 478880 2848
rect 478932 2836 478938 2848
rect 485222 2836 485228 2848
rect 478932 2808 485228 2836
rect 478932 2796 478938 2808
rect 485222 2796 485228 2808
rect 485280 2796 485286 2848
rect 378134 2728 378140 2780
rect 378192 2768 378198 2780
rect 383470 2768 383476 2780
rect 378192 2740 383476 2768
rect 378192 2728 378198 2740
rect 383470 2728 383476 2740
rect 383528 2728 383534 2780
rect 362678 1504 362684 1556
rect 362736 1544 362742 1556
rect 366818 1544 366824 1556
rect 362736 1516 366824 1544
rect 362736 1504 362742 1516
rect 366818 1504 366824 1516
rect 366876 1504 366882 1556
rect 368290 1504 368296 1556
rect 368348 1544 368354 1556
rect 372614 1544 372620 1556
rect 368348 1516 372620 1544
rect 368348 1504 368354 1516
rect 372614 1504 372620 1516
rect 372672 1504 372678 1556
rect 380342 1504 380348 1556
rect 380400 1544 380406 1556
rect 385770 1544 385776 1556
rect 380400 1516 385776 1544
rect 380400 1504 380406 1516
rect 385770 1504 385776 1516
rect 385828 1504 385834 1556
rect 386966 1504 386972 1556
rect 387024 1544 387030 1556
rect 392670 1544 392676 1556
rect 387024 1516 392676 1544
rect 387024 1504 387030 1516
rect 392670 1504 392676 1516
rect 392728 1504 392734 1556
rect 393590 1504 393596 1556
rect 393648 1544 393654 1556
rect 399938 1544 399944 1556
rect 393648 1516 399944 1544
rect 393648 1504 393654 1516
rect 399938 1504 399944 1516
rect 399996 1504 400002 1556
rect 131850 1408 131856 1420
rect 131592 1380 131856 1408
rect 28258 1300 28264 1352
rect 28316 1340 28322 1352
rect 30282 1340 30288 1352
rect 28316 1312 30288 1340
rect 28316 1300 28322 1312
rect 30282 1300 30288 1312
rect 30340 1300 30346 1352
rect 31018 1300 31024 1352
rect 31076 1340 31082 1352
rect 38010 1340 38016 1352
rect 31076 1312 38016 1340
rect 31076 1300 31082 1312
rect 38010 1300 38016 1312
rect 38068 1300 38074 1352
rect 59262 1300 59268 1352
rect 59320 1340 59326 1352
rect 67818 1340 67824 1352
rect 59320 1312 67824 1340
rect 59320 1300 59326 1312
rect 67818 1300 67824 1312
rect 67876 1300 67882 1352
rect 68922 1300 68928 1352
rect 68980 1340 68986 1352
rect 76650 1340 76656 1352
rect 68980 1312 76656 1340
rect 68980 1300 68986 1312
rect 76650 1300 76656 1312
rect 76708 1300 76714 1352
rect 83274 1340 83280 1352
rect 77128 1312 83280 1340
rect 10962 1232 10968 1284
rect 11020 1272 11026 1284
rect 25866 1272 25872 1284
rect 11020 1244 25872 1272
rect 11020 1232 11026 1244
rect 25866 1232 25872 1244
rect 25924 1232 25930 1284
rect 37182 1232 37188 1284
rect 37240 1272 37246 1284
rect 47946 1272 47952 1284
rect 37240 1244 47952 1272
rect 37240 1232 37246 1244
rect 47946 1232 47952 1244
rect 48004 1232 48010 1284
rect 49602 1232 49608 1284
rect 49660 1272 49666 1284
rect 58986 1272 58992 1284
rect 49660 1244 58992 1272
rect 49660 1232 49666 1244
rect 58986 1232 58992 1244
rect 59044 1232 59050 1284
rect 9582 1164 9588 1216
rect 9640 1204 9646 1216
rect 23658 1204 23664 1216
rect 9640 1176 23664 1204
rect 9640 1164 9646 1176
rect 23658 1164 23664 1176
rect 23716 1164 23722 1216
rect 23842 1164 23848 1216
rect 23900 1204 23906 1216
rect 40218 1204 40224 1216
rect 23900 1176 40224 1204
rect 23900 1164 23906 1176
rect 40218 1164 40224 1176
rect 40276 1164 40282 1216
rect 40402 1164 40408 1216
rect 40460 1204 40466 1216
rect 53466 1204 53472 1216
rect 40460 1176 53472 1204
rect 40460 1164 40466 1176
rect 53466 1164 53472 1176
rect 53524 1164 53530 1216
rect 67910 1164 67916 1216
rect 67968 1204 67974 1216
rect 77128 1204 77156 1312
rect 83274 1300 83280 1312
rect 83332 1300 83338 1352
rect 104526 1300 104532 1352
rect 104584 1340 104590 1352
rect 117498 1340 117504 1352
rect 104584 1312 117504 1340
rect 104584 1300 104590 1312
rect 117498 1300 117504 1312
rect 117556 1300 117562 1352
rect 119890 1300 119896 1352
rect 119948 1340 119954 1352
rect 131592 1340 131620 1380
rect 131850 1368 131856 1380
rect 131908 1368 131914 1420
rect 119948 1312 131620 1340
rect 119948 1300 119954 1312
rect 132034 1300 132040 1352
rect 132092 1340 132098 1352
rect 142890 1340 142896 1352
rect 132092 1312 142896 1340
rect 132092 1300 132098 1312
rect 142890 1300 142896 1312
rect 142948 1300 142954 1352
rect 146202 1300 146208 1352
rect 146260 1340 146266 1352
rect 156138 1340 156144 1352
rect 146260 1312 156144 1340
rect 146260 1300 146266 1312
rect 156138 1300 156144 1312
rect 156196 1300 156202 1352
rect 164142 1300 164148 1352
rect 164200 1340 164206 1352
rect 172698 1340 172704 1352
rect 164200 1312 172704 1340
rect 164200 1300 164206 1312
rect 172698 1300 172704 1312
rect 172756 1300 172762 1352
rect 431126 1300 431132 1352
rect 431184 1340 431190 1352
rect 439958 1340 439964 1352
rect 431184 1312 439964 1340
rect 431184 1300 431190 1312
rect 439958 1300 439964 1312
rect 440016 1300 440022 1352
rect 450998 1300 451004 1352
rect 451056 1340 451062 1352
rect 461302 1340 461308 1352
rect 451056 1312 461308 1340
rect 451056 1300 451062 1312
rect 461302 1300 461308 1312
rect 461360 1300 461366 1352
rect 462038 1300 462044 1352
rect 462096 1340 462102 1352
rect 462096 1312 466316 1340
rect 462096 1300 462102 1312
rect 77202 1232 77208 1284
rect 77260 1272 77266 1284
rect 85482 1272 85488 1284
rect 77260 1244 85488 1272
rect 77260 1232 77266 1244
rect 85482 1232 85488 1244
rect 85540 1232 85546 1284
rect 107194 1232 107200 1284
rect 107252 1272 107258 1284
rect 119706 1272 119712 1284
rect 107252 1244 119712 1272
rect 107252 1232 107258 1244
rect 119706 1232 119712 1244
rect 119764 1232 119770 1284
rect 121362 1232 121368 1284
rect 121420 1272 121426 1284
rect 132954 1272 132960 1284
rect 121420 1244 132960 1272
rect 121420 1232 121426 1244
rect 132954 1232 132960 1244
rect 133012 1232 133018 1284
rect 454310 1232 454316 1284
rect 454368 1272 454374 1284
rect 465074 1272 465080 1284
rect 454368 1244 465080 1272
rect 454368 1232 454374 1244
rect 465074 1232 465080 1244
rect 465132 1232 465138 1284
rect 466288 1272 466316 1312
rect 467558 1300 467564 1352
rect 467616 1340 467622 1352
rect 472986 1340 472992 1352
rect 467616 1312 472992 1340
rect 467616 1300 467622 1312
rect 472986 1300 472992 1312
rect 473044 1300 473050 1352
rect 473078 1300 473084 1352
rect 473136 1340 473142 1352
rect 478874 1340 478880 1352
rect 473136 1312 478880 1340
rect 473136 1300 473142 1312
rect 478874 1300 478880 1312
rect 478932 1300 478938 1352
rect 479702 1300 479708 1352
rect 479760 1340 479766 1352
rect 492030 1340 492036 1352
rect 479760 1312 492036 1340
rect 479760 1300 479766 1312
rect 492030 1300 492036 1312
rect 492088 1300 492094 1352
rect 496262 1300 496268 1352
rect 496320 1340 496326 1352
rect 509602 1340 509608 1352
rect 496320 1312 509608 1340
rect 496320 1300 496326 1312
rect 509602 1300 509608 1312
rect 509660 1300 509666 1352
rect 533798 1300 533804 1352
rect 533856 1340 533862 1352
rect 550082 1340 550088 1352
rect 533856 1312 550088 1340
rect 533856 1300 533862 1312
rect 550082 1300 550088 1312
rect 550140 1300 550146 1352
rect 553670 1300 553676 1352
rect 553728 1340 553734 1352
rect 571058 1340 571064 1352
rect 553728 1312 571064 1340
rect 553728 1300 553734 1312
rect 571058 1300 571064 1312
rect 571116 1300 571122 1352
rect 473354 1272 473360 1284
rect 466288 1244 473360 1272
rect 473354 1232 473360 1244
rect 473412 1232 473418 1284
rect 488442 1232 488448 1284
rect 488500 1272 488506 1284
rect 501690 1272 501696 1284
rect 488500 1244 501696 1272
rect 488500 1232 488506 1244
rect 501690 1232 501696 1244
rect 501748 1232 501754 1284
rect 516042 1232 516048 1284
rect 516100 1272 516106 1284
rect 531314 1272 531320 1284
rect 516100 1244 531320 1272
rect 516100 1232 516106 1244
rect 531314 1232 531320 1244
rect 531372 1232 531378 1284
rect 537110 1232 537116 1284
rect 537168 1272 537174 1284
rect 537168 1244 547874 1272
rect 537168 1232 537174 1244
rect 67968 1176 77156 1204
rect 67968 1164 67974 1176
rect 81434 1164 81440 1216
rect 81492 1204 81498 1216
rect 95418 1204 95424 1216
rect 81492 1176 95424 1204
rect 81492 1164 81498 1176
rect 95418 1164 95424 1176
rect 95476 1164 95482 1216
rect 97902 1164 97908 1216
rect 97960 1204 97966 1216
rect 110874 1204 110880 1216
rect 97960 1176 110880 1204
rect 97960 1164 97966 1176
rect 110874 1164 110880 1176
rect 110932 1164 110938 1216
rect 116486 1164 116492 1216
rect 116544 1204 116550 1216
rect 128538 1204 128544 1216
rect 116544 1176 128544 1204
rect 116544 1164 116550 1176
rect 128538 1164 128544 1176
rect 128596 1164 128602 1216
rect 136266 1204 136272 1216
rect 132466 1176 136272 1204
rect 11698 1096 11704 1148
rect 11756 1136 11762 1148
rect 24762 1136 24768 1148
rect 11756 1108 24768 1136
rect 11756 1096 11762 1108
rect 24762 1096 24768 1108
rect 24820 1096 24826 1148
rect 30282 1096 30288 1148
rect 30340 1136 30346 1148
rect 42426 1136 42432 1148
rect 30340 1108 42432 1136
rect 30340 1096 30346 1108
rect 42426 1096 42432 1108
rect 42484 1096 42490 1148
rect 110966 1096 110972 1148
rect 111024 1136 111030 1148
rect 123018 1136 123024 1148
rect 111024 1108 123024 1136
rect 111024 1096 111030 1108
rect 123018 1096 123024 1108
rect 123076 1096 123082 1148
rect 125134 1096 125140 1148
rect 125192 1136 125198 1148
rect 132466 1136 132494 1176
rect 136266 1164 136272 1176
rect 136324 1164 136330 1216
rect 466362 1164 466368 1216
rect 466420 1204 466426 1216
rect 477862 1204 477868 1216
rect 466420 1176 477868 1204
rect 466420 1164 466426 1176
rect 477862 1164 477868 1176
rect 477920 1164 477926 1216
rect 530486 1164 530492 1216
rect 530544 1204 530550 1216
rect 546494 1204 546500 1216
rect 530544 1176 546500 1204
rect 530544 1164 530550 1176
rect 546494 1164 546500 1176
rect 546552 1164 546558 1216
rect 547846 1204 547874 1244
rect 550358 1232 550364 1284
rect 550416 1272 550422 1284
rect 567562 1272 567568 1284
rect 550416 1244 567568 1272
rect 550416 1232 550422 1244
rect 567562 1232 567568 1244
rect 567620 1232 567626 1284
rect 553762 1204 553768 1216
rect 547846 1176 553768 1204
rect 553762 1164 553768 1176
rect 553820 1164 553826 1216
rect 555878 1164 555884 1216
rect 555936 1204 555942 1216
rect 573358 1204 573364 1216
rect 555936 1176 573364 1204
rect 555936 1164 555942 1176
rect 573358 1164 573364 1176
rect 573416 1164 573422 1216
rect 125192 1108 132494 1136
rect 125192 1096 125198 1108
rect 472986 1096 472992 1148
rect 473044 1136 473050 1148
rect 478874 1136 478880 1148
rect 473044 1108 478880 1136
rect 473044 1096 473050 1108
rect 478874 1096 478880 1108
rect 478932 1096 478938 1148
rect 521562 1096 521568 1148
rect 521620 1136 521626 1148
rect 537018 1136 537024 1148
rect 521620 1108 537024 1136
rect 521620 1096 521626 1108
rect 537018 1096 537024 1108
rect 537076 1096 537082 1148
rect 549162 1096 549168 1148
rect 549220 1136 549226 1148
rect 566826 1136 566832 1148
rect 549220 1108 566832 1136
rect 549220 1096 549226 1108
rect 566826 1096 566832 1108
rect 566884 1096 566890 1148
rect 19242 1028 19248 1080
rect 19300 1068 19306 1080
rect 31386 1068 31392 1080
rect 19300 1040 31392 1068
rect 19300 1028 19306 1040
rect 31386 1028 31392 1040
rect 31444 1028 31450 1080
rect 36998 1028 37004 1080
rect 37056 1068 37062 1080
rect 45738 1068 45744 1080
rect 37056 1040 45744 1068
rect 37056 1028 37062 1040
rect 45738 1028 45744 1040
rect 45796 1028 45802 1080
rect 17862 960 17868 1012
rect 17920 1000 17926 1012
rect 28074 1000 28080 1012
rect 17920 972 28080 1000
rect 17920 960 17926 972
rect 28074 960 28080 972
rect 28132 960 28138 1012
rect 33226 960 33232 1012
rect 33284 1000 33290 1012
rect 49050 1000 49056 1012
rect 33284 972 49056 1000
rect 33284 960 33290 972
rect 49050 960 49056 972
rect 49108 960 49114 1012
rect 25774 892 25780 944
rect 25832 932 25838 944
rect 43530 932 43536 944
rect 25832 904 43536 932
rect 25832 892 25838 904
rect 43530 892 43536 904
rect 43588 892 43594 944
rect 9950 824 9956 876
rect 10008 864 10014 876
rect 29178 864 29184 876
rect 10008 836 29184 864
rect 10008 824 10014 836
rect 29178 824 29184 836
rect 29236 824 29242 876
rect 500678 756 500684 808
rect 500736 796 500742 808
rect 514754 796 514760 808
rect 500736 768 514760 796
rect 500736 756 500742 768
rect 514754 756 514760 768
rect 514812 756 514818 808
rect 50154 688 50160 740
rect 50212 728 50218 740
rect 66714 728 66720 740
rect 50212 700 66720 728
rect 50212 688 50218 700
rect 66714 688 66720 700
rect 66772 688 66778 740
rect 497366 688 497372 740
rect 497424 728 497430 740
rect 497424 700 504404 728
rect 497424 688 497430 700
rect 46658 620 46664 672
rect 46716 660 46722 672
rect 63402 660 63408 672
rect 46716 632 63408 660
rect 46716 620 46722 632
rect 63402 620 63408 632
rect 63460 620 63466 672
rect 98638 620 98644 672
rect 98696 660 98702 672
rect 111978 660 111984 672
rect 98696 632 111984 660
rect 98696 620 98702 632
rect 111978 620 111984 632
rect 112036 620 112042 672
rect 482922 620 482928 672
rect 482980 660 482986 672
rect 495894 660 495900 672
rect 482980 632 495900 660
rect 482980 620 482986 632
rect 495894 620 495900 632
rect 495952 620 495958 672
rect 499482 620 499488 672
rect 499540 660 499546 672
rect 499540 620 499574 660
rect 45462 552 45468 604
rect 45520 592 45526 604
rect 62298 592 62304 604
rect 45520 564 62304 592
rect 45520 552 45526 564
rect 62298 552 62304 564
rect 62356 552 62362 604
rect 64322 552 64328 604
rect 64380 592 64386 604
rect 79962 592 79968 604
rect 64380 564 79968 592
rect 64380 552 64386 564
rect 79962 552 79968 564
rect 80020 552 80026 604
rect 99926 552 99932 604
rect 99984 552 99990 604
rect 42886 484 42892 536
rect 42944 524 42950 536
rect 60090 524 60096 536
rect 42944 496 60096 524
rect 42944 484 42950 496
rect 60090 484 60096 496
rect 60148 484 60154 536
rect 63402 484 63408 536
rect 63460 524 63466 536
rect 78858 524 78864 536
rect 63460 496 78864 524
rect 63460 484 63466 496
rect 78858 484 78864 496
rect 78916 484 78922 536
rect 32214 416 32220 468
rect 32272 456 32278 468
rect 49970 456 49976 468
rect 32272 428 49976 456
rect 32272 416 32278 428
rect 49970 416 49976 428
rect 50028 416 50034 468
rect 61838 416 61844 468
rect 61896 456 61902 468
rect 77754 456 77760 468
rect 61896 428 77760 456
rect 61896 416 61902 428
rect 77754 416 77760 428
rect 77812 416 77818 468
rect 86126 416 86132 468
rect 86184 456 86190 468
rect 99944 456 99972 552
rect 86184 428 99972 456
rect 86184 416 86190 428
rect 28718 348 28724 400
rect 28776 388 28782 400
rect 46842 388 46848 400
rect 28776 360 46848 388
rect 28776 348 28782 360
rect 46842 348 46848 360
rect 46900 348 46906 400
rect 48774 348 48780 400
rect 48832 388 48838 400
rect 65702 388 65708 400
rect 48832 360 65708 388
rect 48832 348 48838 360
rect 65702 348 65708 360
rect 65760 348 65766 400
rect 78398 348 78404 400
rect 78456 388 78462 400
rect 93210 388 93216 400
rect 78456 360 93216 388
rect 78456 348 78462 360
rect 93210 348 93216 360
rect 93268 348 93274 400
rect 96062 348 96068 400
rect 96120 388 96126 400
rect 109770 388 109776 400
rect 96120 360 109776 388
rect 96120 348 96126 360
rect 109770 348 109776 360
rect 109828 348 109834 400
rect 20438 280 20444 332
rect 20496 320 20502 332
rect 39114 320 39120 332
rect 20496 292 39120 320
rect 20496 280 20502 292
rect 39114 280 39120 292
rect 39172 280 39178 332
rect 39390 280 39396 332
rect 39448 320 39454 332
rect 56778 320 56784 332
rect 39448 292 56784 320
rect 39448 280 39454 292
rect 56778 280 56784 292
rect 56836 280 56842 332
rect 57054 280 57060 332
rect 57112 320 57118 332
rect 73338 320 73344 332
rect 57112 292 73344 320
rect 57112 280 57118 292
rect 73338 280 73344 292
rect 73396 280 73402 332
rect 79502 280 79508 332
rect 79560 320 79566 332
rect 94314 320 94320 332
rect 79560 292 94320 320
rect 79560 280 79566 292
rect 94314 280 94320 292
rect 94372 280 94378 332
rect 94958 280 94964 332
rect 95016 320 95022 332
rect 108666 320 108672 332
rect 95016 292 108672 320
rect 95016 280 95022 292
rect 108666 280 108672 292
rect 108724 280 108730 332
rect 499546 320 499574 620
rect 504376 456 504404 700
rect 513926 688 513932 740
rect 513984 728 513990 740
rect 529014 728 529020 740
rect 513984 700 529020 728
rect 513984 688 513990 700
rect 529014 688 529020 700
rect 529072 688 529078 740
rect 520734 660 520740 672
rect 518866 632 520740 660
rect 511442 456 511448 468
rect 504376 428 511448 456
rect 511442 416 511448 428
rect 511500 416 511506 468
rect 506198 348 506204 400
rect 506256 388 506262 400
rect 518866 388 518894 632
rect 520734 620 520740 632
rect 520792 620 520798 672
rect 539318 416 539324 468
rect 539376 456 539382 468
rect 556338 456 556344 468
rect 539376 428 556344 456
rect 539376 416 539382 428
rect 556338 416 556344 428
rect 556396 416 556402 468
rect 506256 360 518894 388
rect 506256 348 506262 360
rect 523862 348 523868 400
rect 523920 388 523926 400
rect 539778 388 539784 400
rect 523920 360 539784 388
rect 523920 348 523926 360
rect 539778 348 539784 360
rect 539836 348 539842 400
rect 547046 348 547052 400
rect 547104 388 547110 400
rect 564618 388 564624 400
rect 547104 360 564624 388
rect 547104 348 547110 360
rect 564618 348 564624 360
rect 564676 348 564682 400
rect 513374 320 513380 332
rect 499546 292 513380 320
rect 513374 280 513380 292
rect 513432 280 513438 332
rect 517330 280 517336 332
rect 517388 320 517394 332
rect 532142 320 532148 332
rect 517388 292 532148 320
rect 517388 280 517394 292
rect 532142 280 532148 292
rect 532200 280 532206 332
rect 532694 280 532700 332
rect 532752 320 532758 332
rect 548702 320 548708 332
rect 532752 292 548708 320
rect 532752 280 532758 292
rect 548702 280 548708 292
rect 548760 280 548766 332
rect 554682 280 554688 332
rect 554740 320 554746 332
rect 572898 320 572904 332
rect 554740 292 572904 320
rect 554740 280 554746 292
rect 572898 280 572904 292
rect 572956 280 572962 332
rect 16206 212 16212 264
rect 16264 252 16270 264
rect 34606 252 34612 264
rect 16264 224 34612 252
rect 16264 212 16270 224
rect 34606 212 34612 224
rect 34664 212 34670 264
rect 38562 212 38568 264
rect 38620 252 38626 264
rect 55674 252 55680 264
rect 38620 224 55680 252
rect 38620 212 38626 224
rect 55674 212 55680 224
rect 55732 212 55738 264
rect 56410 212 56416 264
rect 56468 252 56474 264
rect 72234 252 72240 264
rect 56468 224 72240 252
rect 56468 212 56474 224
rect 72234 212 72240 224
rect 72292 212 72298 264
rect 75362 212 75368 264
rect 75420 252 75426 264
rect 89898 252 89904 264
rect 75420 224 89904 252
rect 75420 212 75426 224
rect 89898 212 89904 224
rect 89956 212 89962 264
rect 92566 212 92572 264
rect 92624 252 92630 264
rect 106458 252 106464 264
rect 92624 224 106464 252
rect 92624 212 92630 224
rect 106458 212 106464 224
rect 106516 212 106522 264
rect 484210 212 484216 264
rect 484268 252 484274 264
rect 497274 252 497280 264
rect 484268 224 497280 252
rect 484268 212 484274 224
rect 497274 212 497280 224
rect 497332 212 497338 264
rect 505002 212 505008 264
rect 505060 252 505066 264
rect 519722 252 519728 264
rect 505060 224 519728 252
rect 505060 212 505066 224
rect 519722 212 519728 224
rect 519780 212 519786 264
rect 520550 212 520556 264
rect 520608 252 520614 264
rect 536282 252 536288 264
rect 520608 224 536288 252
rect 520608 212 520614 224
rect 536282 212 536288 224
rect 536340 212 536346 264
rect 538122 212 538128 264
rect 538180 252 538186 264
rect 554774 252 554780 264
rect 538180 224 554780 252
rect 538180 212 538186 224
rect 554774 212 554780 224
rect 554832 212 554838 264
rect 556890 212 556896 264
rect 556948 252 556954 264
rect 575290 252 575296 264
rect 556948 224 575296 252
rect 556948 212 556954 224
rect 575290 212 575296 224
rect 575348 212 575354 264
rect 14550 144 14556 196
rect 14608 184 14614 196
rect 33410 184 33416 196
rect 14608 156 33416 184
rect 14608 144 14614 156
rect 33410 144 33416 156
rect 33468 144 33474 196
rect 36998 144 37004 196
rect 37056 184 37062 196
rect 54570 184 54576 196
rect 37056 156 54576 184
rect 37056 144 37062 156
rect 54570 144 54576 156
rect 54628 144 54634 196
rect 55122 144 55128 196
rect 55180 184 55186 196
rect 71130 184 71136 196
rect 55180 156 71136 184
rect 55180 144 55186 156
rect 71130 144 71136 156
rect 71188 144 71194 196
rect 73614 144 73620 196
rect 73672 184 73678 196
rect 88794 184 88800 196
rect 73672 156 88800 184
rect 73672 144 73678 156
rect 88794 144 88800 156
rect 88852 144 88858 196
rect 89530 144 89536 196
rect 89588 184 89594 196
rect 103146 184 103152 196
rect 89588 156 103152 184
rect 89588 144 89594 156
rect 103146 144 103152 156
rect 103204 144 103210 196
rect 114370 144 114376 196
rect 114428 184 114434 196
rect 126330 184 126336 196
rect 114428 156 126336 184
rect 114428 144 114434 156
rect 126330 144 126336 156
rect 126388 144 126394 196
rect 128354 144 128360 196
rect 128412 184 128418 196
rect 139578 184 139584 196
rect 128412 156 139584 184
rect 128412 144 128418 156
rect 139578 144 139584 156
rect 139636 144 139642 196
rect 144914 144 144920 196
rect 144972 184 144978 196
rect 155034 184 155040 196
rect 144972 156 155040 184
rect 144972 144 144978 156
rect 155034 144 155040 156
rect 155092 144 155098 196
rect 438762 144 438768 196
rect 438820 184 438826 196
rect 448422 184 448428 196
rect 438820 156 448428 184
rect 438820 144 438826 156
rect 448422 144 448428 156
rect 448480 144 448486 196
rect 474182 144 474188 196
rect 474240 184 474246 196
rect 486602 184 486608 196
rect 474240 156 486608 184
rect 474240 144 474246 156
rect 486602 144 486608 156
rect 486660 144 486666 196
rect 490650 144 490656 196
rect 490708 184 490714 196
rect 503806 184 503812 196
rect 490708 156 503812 184
rect 490708 144 490714 156
rect 503806 144 503812 156
rect 503864 144 503870 196
rect 507210 144 507216 196
rect 507268 184 507274 196
rect 521654 184 521660 196
rect 507268 156 521660 184
rect 507268 144 507274 156
rect 521654 144 521660 156
rect 521712 144 521718 196
rect 522758 144 522764 196
rect 522816 184 522822 196
rect 538214 184 538220 196
rect 522816 156 538220 184
rect 522816 144 522822 156
rect 538214 144 538220 156
rect 538272 144 538278 196
rect 540422 144 540428 196
rect 540480 184 540486 196
rect 556982 184 556988 196
rect 540480 156 556988 184
rect 540480 144 540486 156
rect 556982 144 556988 156
rect 557040 144 557046 196
rect 560202 144 560208 196
rect 560260 184 560266 196
rect 578786 184 578792 196
rect 560260 156 578792 184
rect 560260 144 560266 156
rect 578786 144 578792 156
rect 578844 144 578850 196
rect 13722 76 13728 128
rect 13780 116 13786 128
rect 32582 116 32588 128
rect 13780 88 32588 116
rect 13780 76 13786 88
rect 32582 76 32588 88
rect 32640 76 32646 128
rect 33778 76 33784 128
rect 33836 116 33842 128
rect 51166 116 51172 128
rect 33836 88 51172 116
rect 33836 76 33842 88
rect 51166 76 51172 88
rect 51224 76 51230 128
rect 53558 76 53564 128
rect 53616 116 53622 128
rect 70026 116 70032 128
rect 53616 88 70032 116
rect 53616 76 53622 88
rect 70026 76 70032 88
rect 70084 76 70090 128
rect 71682 76 71688 128
rect 71740 116 71746 128
rect 86586 116 86592 128
rect 71740 88 86592 116
rect 71740 76 71746 88
rect 86586 76 86592 88
rect 86644 76 86650 128
rect 86678 76 86684 128
rect 86736 116 86742 128
rect 100846 116 100852 128
rect 86736 88 100852 116
rect 86736 76 86742 88
rect 100846 76 100852 88
rect 100904 76 100910 128
rect 103514 76 103520 128
rect 103572 116 103578 128
rect 116210 116 116216 128
rect 103572 88 116216 116
rect 103572 76 103578 88
rect 116210 76 116216 88
rect 116268 76 116274 128
rect 122558 76 122564 128
rect 122616 116 122622 128
rect 133966 116 133972 128
rect 122616 88 133972 116
rect 122616 76 122622 88
rect 133966 76 133972 88
rect 134024 76 134030 128
rect 139210 76 139216 128
rect 139268 116 139274 128
rect 149330 116 149336 128
rect 139268 88 149336 116
rect 139268 76 139274 88
rect 149330 76 149336 88
rect 149388 76 149394 128
rect 422202 76 422208 128
rect 422260 116 422266 128
rect 431034 116 431040 128
rect 422260 88 431040 116
rect 422260 76 422266 88
rect 431034 76 431040 88
rect 431092 76 431098 128
rect 444282 76 444288 128
rect 444340 116 444346 128
rect 454126 116 454132 128
rect 444340 88 454132 116
rect 444340 76 444346 88
rect 454126 76 454132 88
rect 454184 76 454190 128
rect 460842 76 460848 128
rect 460900 116 460906 128
rect 472434 116 472440 128
rect 460900 88 472440 116
rect 460900 76 460906 88
rect 472434 76 472440 88
rect 472492 76 472498 128
rect 477402 76 477408 128
rect 477460 116 477466 128
rect 490098 116 490104 128
rect 477460 88 490104 116
rect 477460 76 477466 88
rect 490098 76 490104 88
rect 490156 76 490162 128
rect 493962 76 493968 128
rect 494020 116 494026 128
rect 507302 116 507308 128
rect 494020 88 507308 116
rect 494020 76 494026 88
rect 507302 76 507308 88
rect 507360 76 507366 128
rect 510522 76 510528 128
rect 510580 116 510586 128
rect 525610 116 525616 128
rect 510580 88 525616 116
rect 510580 76 510586 88
rect 525610 76 525616 88
rect 525668 76 525674 128
rect 527082 76 527088 128
rect 527140 116 527146 128
rect 542814 116 542820 128
rect 527140 88 542820 116
rect 527140 76 527146 88
rect 542814 76 542820 88
rect 542872 76 542878 128
rect 543642 76 543648 128
rect 543700 116 543706 128
rect 560478 116 560484 128
rect 543700 88 560484 116
rect 543700 76 543706 88
rect 560478 76 560484 88
rect 560536 76 560542 128
rect 561398 76 561404 128
rect 561456 116 561462 128
rect 581178 116 581184 128
rect 561456 88 581184 116
rect 561456 76 561462 88
rect 581178 76 581184 88
rect 581236 76 581242 128
<< via1 >>
rect 35992 2864 36044 2916
rect 40408 2864 40460 2916
rect 134340 2864 134392 2916
rect 145150 2864 145202 2916
rect 169576 2864 169628 2916
rect 178270 2864 178322 2916
rect 359326 2864 359378 2916
rect 363328 2864 363380 2916
rect 364064 2864 364116 2916
rect 365720 2864 365772 2916
rect 365950 2864 366002 2916
rect 370044 2864 370096 2916
rect 370366 2864 370418 2916
rect 375196 2864 375248 2916
rect 376990 2864 377042 2916
rect 382280 2864 382332 2916
rect 385822 2864 385874 2916
rect 391848 2864 391900 2916
rect 393228 2864 393280 2916
rect 394056 2864 394108 2916
rect 394654 2864 394706 2916
rect 400864 2864 400916 2916
rect 30104 2796 30156 2848
rect 37188 2796 37240 2848
rect 41880 2796 41932 2848
rect 49608 2796 49660 2848
rect 51356 2796 51408 2848
rect 59268 2796 59320 2848
rect 60832 2796 60884 2848
rect 68928 2796 68980 2848
rect 70308 2796 70360 2848
rect 77208 2796 77260 2848
rect 82084 2796 82136 2848
rect 96574 2796 96626 2848
rect 153016 2796 153068 2848
rect 162814 2796 162866 2848
rect 351598 2796 351650 2848
rect 355048 2796 355100 2848
rect 358222 2796 358274 2848
rect 361672 2796 361724 2848
rect 367054 2796 367106 2848
rect 371240 2796 371292 2848
rect 371332 2796 371384 2848
rect 374000 2796 374052 2848
rect 375886 2796 375938 2848
rect 380900 2796 380952 2848
rect 389134 2796 389186 2848
rect 393504 2796 393556 2848
rect 395758 2796 395810 2848
rect 402336 2796 402388 2848
rect 404590 2796 404642 2848
rect 411720 2796 411772 2848
rect 449854 2796 449906 2848
rect 460388 2796 460440 2848
rect 478880 2796 478932 2848
rect 485228 2796 485280 2848
rect 378140 2728 378192 2780
rect 383476 2728 383528 2780
rect 362684 1504 362736 1556
rect 366824 1504 366876 1556
rect 368296 1504 368348 1556
rect 372620 1504 372672 1556
rect 380348 1504 380400 1556
rect 385776 1504 385828 1556
rect 386972 1504 387024 1556
rect 392676 1504 392728 1556
rect 393596 1504 393648 1556
rect 399944 1504 399996 1556
rect 28264 1300 28316 1352
rect 30288 1300 30340 1352
rect 31024 1300 31076 1352
rect 38016 1300 38068 1352
rect 59268 1300 59320 1352
rect 67824 1300 67876 1352
rect 68928 1300 68980 1352
rect 76656 1300 76708 1352
rect 10968 1232 11020 1284
rect 25872 1232 25924 1284
rect 37188 1232 37240 1284
rect 47952 1232 48004 1284
rect 49608 1232 49660 1284
rect 58992 1232 59044 1284
rect 9588 1164 9640 1216
rect 23664 1164 23716 1216
rect 23848 1164 23900 1216
rect 40224 1164 40276 1216
rect 40408 1164 40460 1216
rect 53472 1164 53524 1216
rect 67916 1164 67968 1216
rect 83280 1300 83332 1352
rect 104532 1300 104584 1352
rect 117504 1300 117556 1352
rect 119896 1300 119948 1352
rect 131856 1368 131908 1420
rect 132040 1300 132092 1352
rect 142896 1300 142948 1352
rect 146208 1300 146260 1352
rect 156144 1300 156196 1352
rect 164148 1300 164200 1352
rect 172704 1300 172756 1352
rect 431132 1300 431184 1352
rect 439964 1300 440016 1352
rect 451004 1300 451056 1352
rect 461308 1300 461360 1352
rect 462044 1300 462096 1352
rect 77208 1232 77260 1284
rect 85488 1232 85540 1284
rect 107200 1232 107252 1284
rect 119712 1232 119764 1284
rect 121368 1232 121420 1284
rect 132960 1232 133012 1284
rect 454316 1232 454368 1284
rect 465080 1232 465132 1284
rect 467564 1300 467616 1352
rect 472992 1300 473044 1352
rect 473084 1300 473136 1352
rect 478880 1300 478932 1352
rect 479708 1300 479760 1352
rect 492036 1300 492088 1352
rect 496268 1300 496320 1352
rect 509608 1300 509660 1352
rect 533804 1300 533856 1352
rect 550088 1300 550140 1352
rect 553676 1300 553728 1352
rect 571064 1300 571116 1352
rect 473360 1232 473412 1284
rect 488448 1232 488500 1284
rect 501696 1232 501748 1284
rect 516048 1232 516100 1284
rect 531320 1232 531372 1284
rect 537116 1232 537168 1284
rect 81440 1164 81492 1216
rect 95424 1164 95476 1216
rect 97908 1164 97960 1216
rect 110880 1164 110932 1216
rect 116492 1164 116544 1216
rect 128544 1164 128596 1216
rect 11704 1096 11756 1148
rect 24768 1096 24820 1148
rect 30288 1096 30340 1148
rect 42432 1096 42484 1148
rect 110972 1096 111024 1148
rect 123024 1096 123076 1148
rect 125140 1096 125192 1148
rect 136272 1164 136324 1216
rect 466368 1164 466420 1216
rect 477868 1164 477920 1216
rect 530492 1164 530544 1216
rect 546500 1164 546552 1216
rect 550364 1232 550416 1284
rect 567568 1232 567620 1284
rect 553768 1164 553820 1216
rect 555884 1164 555936 1216
rect 573364 1164 573416 1216
rect 472992 1096 473044 1148
rect 478880 1096 478932 1148
rect 521568 1096 521620 1148
rect 537024 1096 537076 1148
rect 549168 1096 549220 1148
rect 566832 1096 566884 1148
rect 19248 1028 19300 1080
rect 31392 1028 31444 1080
rect 37004 1028 37056 1080
rect 45744 1028 45796 1080
rect 17868 960 17920 1012
rect 28080 960 28132 1012
rect 33232 960 33284 1012
rect 49056 960 49108 1012
rect 25780 892 25832 944
rect 43536 892 43588 944
rect 9956 824 10008 876
rect 29184 824 29236 876
rect 500684 756 500736 808
rect 514760 756 514812 808
rect 50160 688 50212 740
rect 66720 688 66772 740
rect 497372 688 497424 740
rect 46664 620 46716 672
rect 63408 620 63460 672
rect 98644 620 98696 672
rect 111984 620 112036 672
rect 482928 620 482980 672
rect 495900 620 495952 672
rect 499488 620 499540 672
rect 45468 552 45520 604
rect 62304 552 62356 604
rect 64328 552 64380 604
rect 79968 552 80020 604
rect 99932 552 99984 604
rect 42892 484 42944 536
rect 60096 484 60148 536
rect 63408 484 63460 536
rect 78864 484 78916 536
rect 32220 416 32272 468
rect 49976 416 50028 468
rect 61844 416 61896 468
rect 77760 416 77812 468
rect 86132 416 86184 468
rect 28724 348 28776 400
rect 46848 348 46900 400
rect 48780 348 48832 400
rect 65708 348 65760 400
rect 78404 348 78456 400
rect 93216 348 93268 400
rect 96068 348 96120 400
rect 109776 348 109828 400
rect 20444 280 20496 332
rect 39120 280 39172 332
rect 39396 280 39448 332
rect 56784 280 56836 332
rect 57060 280 57112 332
rect 73344 280 73396 332
rect 79508 280 79560 332
rect 94320 280 94372 332
rect 94964 280 95016 332
rect 108672 280 108724 332
rect 513932 688 513984 740
rect 529020 688 529072 740
rect 511448 416 511500 468
rect 506204 348 506256 400
rect 520740 620 520792 672
rect 539324 416 539376 468
rect 556344 416 556396 468
rect 523868 348 523920 400
rect 539784 348 539836 400
rect 547052 348 547104 400
rect 564624 348 564676 400
rect 513380 280 513432 332
rect 517336 280 517388 332
rect 532148 280 532200 332
rect 532700 280 532752 332
rect 548708 280 548760 332
rect 554688 280 554740 332
rect 572904 280 572956 332
rect 16212 212 16264 264
rect 34612 212 34664 264
rect 38568 212 38620 264
rect 55680 212 55732 264
rect 56416 212 56468 264
rect 72240 212 72292 264
rect 75368 212 75420 264
rect 89904 212 89956 264
rect 92572 212 92624 264
rect 106464 212 106516 264
rect 484216 212 484268 264
rect 497280 212 497332 264
rect 505008 212 505060 264
rect 519728 212 519780 264
rect 520556 212 520608 264
rect 536288 212 536340 264
rect 538128 212 538180 264
rect 554780 212 554832 264
rect 556896 212 556948 264
rect 575296 212 575348 264
rect 14556 144 14608 196
rect 33416 144 33468 196
rect 37004 144 37056 196
rect 54576 144 54628 196
rect 55128 144 55180 196
rect 71136 144 71188 196
rect 73620 144 73672 196
rect 88800 144 88852 196
rect 89536 144 89588 196
rect 103152 144 103204 196
rect 114376 144 114428 196
rect 126336 144 126388 196
rect 128360 144 128412 196
rect 139584 144 139636 196
rect 144920 144 144972 196
rect 155040 144 155092 196
rect 438768 144 438820 196
rect 448428 144 448480 196
rect 474188 144 474240 196
rect 486608 144 486660 196
rect 490656 144 490708 196
rect 503812 144 503864 196
rect 507216 144 507268 196
rect 521660 144 521712 196
rect 522764 144 522816 196
rect 538220 144 538272 196
rect 540428 144 540480 196
rect 556988 144 557040 196
rect 560208 144 560260 196
rect 578792 144 578844 196
rect 13728 76 13780 128
rect 32588 76 32640 128
rect 33784 76 33836 128
rect 51172 76 51224 128
rect 53564 76 53616 128
rect 70032 76 70084 128
rect 71688 76 71740 128
rect 86592 76 86644 128
rect 86684 76 86736 128
rect 100852 76 100904 128
rect 103520 76 103572 128
rect 116216 76 116268 128
rect 122564 76 122616 128
rect 133972 76 134024 128
rect 139216 76 139268 128
rect 149336 76 149388 128
rect 422208 76 422260 128
rect 431040 76 431092 128
rect 444288 76 444340 128
rect 454132 76 454184 128
rect 460848 76 460900 128
rect 472440 76 472492 128
rect 477408 76 477460 128
rect 490104 76 490156 128
rect 493968 76 494020 128
rect 507308 76 507360 128
rect 510528 76 510580 128
rect 525616 76 525668 128
rect 527088 76 527140 128
rect 542820 76 542872 128
rect 543648 76 543700 128
rect 560484 76 560536 128
rect 561404 76 561456 128
rect 581184 76 581236 128
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 17038 2816 17094 2825
rect 20410 2802 20438 3060
rect 21514 2802 21542 3060
rect 22618 2802 22646 3060
rect 17038 2751 17094 2760
rect 20364 2774 20438 2802
rect 21468 2774 21542 2802
rect 22572 2774 22646 2802
rect 23018 2816 23074 2825
rect 10968 1284 11020 1290
rect 10968 1226 11020 1232
rect 9588 1216 9640 1222
rect 9588 1158 9640 1164
rect 6458 1048 6514 1057
rect 6458 983 6514 992
rect 5262 912 5318 921
rect 5262 847 5318 856
rect 4066 640 4122 649
rect 4066 575 4122 584
rect 4080 480 4108 575
rect 5276 480 5304 847
rect 6472 480 6500 983
rect 8758 776 8814 785
rect 8758 711 8814 720
rect 8206 504 8262 513
rect 386 96 442 105
rect 542 82 654 480
rect 1490 232 1546 241
rect 1646 218 1758 480
rect 1546 190 1758 218
rect 1490 167 1546 176
rect 442 54 654 82
rect 386 31 442 40
rect 542 -960 654 54
rect 1646 -960 1758 190
rect 2842 354 2954 480
rect 3330 368 3386 377
rect 2842 326 3330 354
rect 2842 -960 2954 326
rect 3330 303 3386 312
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 354 7738 480
rect 8128 462 8206 490
rect 8128 354 8156 462
rect 8772 480 8800 711
rect 9600 649 9628 1158
rect 10980 1057 11008 1226
rect 11704 1148 11756 1154
rect 11704 1090 11756 1096
rect 10966 1048 11022 1057
rect 10966 983 11022 992
rect 11716 921 11744 1090
rect 12346 1048 12402 1057
rect 12346 983 12402 992
rect 11702 912 11758 921
rect 9956 876 10008 882
rect 11702 847 11758 856
rect 9956 818 10008 824
rect 9586 640 9642 649
rect 9586 575 9642 584
rect 9968 480 9996 818
rect 11150 640 11206 649
rect 11150 575 11206 584
rect 11164 480 11192 575
rect 12360 480 12388 983
rect 17052 480 17080 2751
rect 19248 1080 19300 1086
rect 19246 1048 19248 1057
rect 19300 1048 19302 1057
rect 17868 1012 17920 1018
rect 19246 983 19302 992
rect 17868 954 17920 960
rect 17880 785 17908 954
rect 19430 912 19486 921
rect 19430 847 19486 856
rect 17866 776 17922 785
rect 17866 711 17922 720
rect 18234 776 18290 785
rect 18234 711 18290 720
rect 18248 480 18276 711
rect 19444 480 19472 847
rect 8206 439 8262 448
rect 7626 326 8156 354
rect 7626 -960 7738 326
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 82 13626 480
rect 14710 218 14822 480
rect 14568 202 14822 218
rect 14556 196 14822 202
rect 14608 190 14822 196
rect 14556 138 14608 144
rect 13728 128 13780 134
rect 13514 76 13728 82
rect 13514 70 13780 76
rect 13514 54 13768 70
rect 13514 -960 13626 54
rect 14710 -960 14822 190
rect 15906 218 16018 480
rect 16212 264 16264 270
rect 15906 212 16212 218
rect 15906 206 16264 212
rect 15906 190 16252 206
rect 15906 -960 16018 190
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20364 105 20392 2774
rect 20598 354 20710 480
rect 20456 338 20710 354
rect 20444 332 20710 338
rect 20496 326 20710 332
rect 20444 274 20496 280
rect 20350 96 20406 105
rect 20350 31 20406 40
rect 20598 -960 20710 326
rect 21468 241 21496 2774
rect 21822 1048 21878 1057
rect 21822 983 21878 992
rect 21836 480 21864 983
rect 21454 232 21510 241
rect 21454 167 21510 176
rect 21794 -960 21906 480
rect 22572 377 22600 2774
rect 23722 2802 23750 3060
rect 24826 2802 24854 3060
rect 25930 2802 25958 3060
rect 27034 2802 27062 3060
rect 28138 2802 28166 3060
rect 29242 2802 29270 3060
rect 23018 2751 23074 2760
rect 23676 2774 23750 2802
rect 24780 2774 24854 2802
rect 25884 2774 25958 2802
rect 26988 2774 27062 2802
rect 28092 2774 28166 2802
rect 29196 2774 29270 2802
rect 30104 2848 30156 2854
rect 30346 2802 30374 3060
rect 31450 2802 31478 3060
rect 30104 2790 30156 2796
rect 23032 480 23060 2751
rect 23676 1222 23704 2774
rect 23664 1216 23716 1222
rect 23664 1158 23716 1164
rect 23848 1216 23900 1222
rect 23848 1158 23900 1164
rect 23860 1057 23888 1158
rect 24780 1154 24808 2774
rect 25884 1290 25912 2774
rect 25872 1284 25924 1290
rect 25872 1226 25924 1232
rect 24768 1148 24820 1154
rect 24768 1090 24820 1096
rect 23846 1048 23902 1057
rect 23846 983 23902 992
rect 25780 944 25832 950
rect 25780 886 25832 892
rect 22558 368 22614 377
rect 22558 303 22614 312
rect 22990 -960 23102 480
rect 24186 354 24298 480
rect 24766 368 24822 377
rect 24186 326 24766 354
rect 24186 -960 24298 326
rect 24766 303 24822 312
rect 25290 354 25402 480
rect 25792 354 25820 886
rect 26988 513 27016 2774
rect 28092 1018 28120 2774
rect 28264 1352 28316 1358
rect 28264 1294 28316 1300
rect 28080 1012 28132 1018
rect 28080 954 28132 960
rect 28276 649 28304 1294
rect 29196 882 29224 2774
rect 29184 876 29236 882
rect 29184 818 29236 824
rect 28262 640 28318 649
rect 28262 575 28318 584
rect 26974 504 27030 513
rect 25290 326 25820 354
rect 25290 -960 25402 326
rect 26330 232 26386 241
rect 26486 218 26598 480
rect 28170 504 28226 513
rect 26974 439 27030 448
rect 26386 190 26598 218
rect 26330 167 26386 176
rect 26486 -960 26598 190
rect 27682 354 27794 480
rect 30116 480 30144 2790
rect 30300 2774 30374 2802
rect 31404 2774 31478 2802
rect 32554 2802 32582 3060
rect 33658 2802 33686 3060
rect 34762 2802 34790 3060
rect 35866 2961 35894 3060
rect 35852 2952 35908 2961
rect 35852 2887 35908 2896
rect 35992 2916 36044 2922
rect 35992 2858 36044 2864
rect 32554 2774 32628 2802
rect 30300 1358 30328 2774
rect 30288 1352 30340 1358
rect 30288 1294 30340 1300
rect 31024 1352 31076 1358
rect 31024 1294 31076 1300
rect 30288 1148 30340 1154
rect 30288 1090 30340 1096
rect 28170 439 28226 448
rect 28184 354 28212 439
rect 27682 326 28212 354
rect 28724 400 28776 406
rect 28878 354 28990 480
rect 28776 348 28990 354
rect 28724 342 28990 348
rect 28736 326 28990 342
rect 27682 -960 27794 326
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30300 377 30328 1090
rect 31036 921 31064 1294
rect 31404 1086 31432 2774
rect 31392 1080 31444 1086
rect 31392 1022 31444 1028
rect 31022 912 31078 921
rect 31022 847 31078 856
rect 31298 640 31354 649
rect 31298 575 31354 584
rect 31312 480 31340 575
rect 30286 368 30342 377
rect 30286 303 30342 312
rect 31270 -960 31382 480
rect 32220 468 32272 474
rect 32220 410 32272 416
rect 32232 354 32260 410
rect 32374 354 32486 480
rect 32232 326 32486 354
rect 32374 -960 32486 326
rect 32600 134 32628 2774
rect 33428 2774 33686 2802
rect 34624 2774 34790 2802
rect 33232 1012 33284 1018
rect 33232 954 33284 960
rect 33244 649 33272 954
rect 33230 640 33286 649
rect 33230 575 33286 584
rect 33428 202 33456 2774
rect 33612 598 33824 626
rect 33612 480 33640 598
rect 33416 196 33468 202
rect 33416 138 33468 144
rect 32588 128 32640 134
rect 32588 70 32640 76
rect 33570 -960 33682 480
rect 33796 134 33824 598
rect 34624 270 34652 2774
rect 34794 2544 34850 2553
rect 34794 2479 34850 2488
rect 34808 480 34836 2479
rect 36004 480 36032 2858
rect 36970 2802 36998 3060
rect 36924 2774 36998 2802
rect 37188 2848 37240 2854
rect 38074 2802 38102 3060
rect 39178 2802 39206 3060
rect 40282 2802 40310 3060
rect 40408 2916 40460 2922
rect 40408 2858 40460 2864
rect 37188 2790 37240 2796
rect 36924 785 36952 2774
rect 37200 1290 37228 2790
rect 38028 2774 38102 2802
rect 39132 2774 39206 2802
rect 40236 2774 40310 2802
rect 38028 1358 38056 2774
rect 38016 1352 38068 1358
rect 38016 1294 38068 1300
rect 37188 1284 37240 1290
rect 37188 1226 37240 1232
rect 37004 1080 37056 1086
rect 37004 1022 37056 1028
rect 36910 776 36966 785
rect 36910 711 36966 720
rect 37016 513 37044 1022
rect 37002 504 37058 513
rect 34612 264 34664 270
rect 34612 206 34664 212
rect 33784 128 33836 134
rect 33784 70 33836 76
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37002 439 37058 448
rect 37158 218 37270 480
rect 37016 202 37270 218
rect 37004 196 37270 202
rect 37056 190 37270 196
rect 37004 138 37056 144
rect 37158 -960 37270 190
rect 38354 218 38466 480
rect 39132 338 39160 2774
rect 40236 1222 40264 2774
rect 40420 1222 40448 2858
rect 41386 2825 41414 3060
rect 41880 2848 41932 2854
rect 41372 2816 41428 2825
rect 42490 2802 42518 3060
rect 43594 2802 43622 3060
rect 44698 2802 44726 3060
rect 45802 2802 45830 3060
rect 46906 2802 46934 3060
rect 48010 2802 48038 3060
rect 49114 2802 49142 3060
rect 41880 2790 41932 2796
rect 41372 2751 41428 2760
rect 40774 2680 40830 2689
rect 40696 2638 40774 2666
rect 40224 1216 40276 1222
rect 40224 1158 40276 1164
rect 40408 1216 40460 1222
rect 40408 1158 40460 1164
rect 40696 480 40724 2638
rect 40774 2615 40830 2624
rect 41892 480 41920 2790
rect 42444 2774 42518 2802
rect 43548 2774 43622 2802
rect 44652 2774 44726 2802
rect 45756 2774 45830 2802
rect 46860 2774 46934 2802
rect 47964 2774 48038 2802
rect 49068 2774 49142 2802
rect 49608 2848 49660 2854
rect 50218 2802 50246 3060
rect 51322 2938 51350 3060
rect 52426 2961 52454 3060
rect 49608 2790 49660 2796
rect 42444 1154 42472 2774
rect 42432 1148 42484 1154
rect 42432 1090 42484 1096
rect 43548 950 43576 2774
rect 43536 944 43588 950
rect 43536 886 43588 892
rect 42892 536 42944 542
rect 39550 354 39662 480
rect 39408 338 39662 354
rect 39120 332 39172 338
rect 39120 274 39172 280
rect 39396 332 39662 338
rect 39448 326 39662 332
rect 39396 274 39448 280
rect 38568 264 38620 270
rect 38354 212 38568 218
rect 38354 206 38620 212
rect 38354 190 38608 206
rect 38354 -960 38466 190
rect 39550 -960 39662 326
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 42892 478 42944 484
rect 42904 354 42932 478
rect 43046 354 43158 480
rect 42904 326 43158 354
rect 43046 -960 43158 326
rect 44242 82 44354 480
rect 44652 241 44680 2774
rect 45756 1086 45784 2774
rect 45744 1080 45796 1086
rect 45744 1022 45796 1028
rect 46664 672 46716 678
rect 46664 614 46716 620
rect 45468 604 45520 610
rect 45468 546 45520 552
rect 45480 480 45508 546
rect 46676 480 46704 614
rect 44638 232 44694 241
rect 44638 167 44694 176
rect 44638 96 44694 105
rect 44242 54 44638 82
rect 44242 -960 44354 54
rect 44638 31 44694 40
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 46860 406 46888 2774
rect 47858 2680 47914 2689
rect 47858 2615 47914 2624
rect 47872 480 47900 2615
rect 47964 1290 47992 2774
rect 47952 1284 48004 1290
rect 47952 1226 48004 1232
rect 49068 1018 49096 2774
rect 49620 1290 49648 2790
rect 49988 2774 50246 2802
rect 51184 2910 51350 2938
rect 52412 2952 52468 2961
rect 49608 1284 49660 1290
rect 49608 1226 49660 1232
rect 49056 1012 49108 1018
rect 49056 954 49108 960
rect 46848 400 46900 406
rect 46848 342 46900 348
rect 47830 -960 47942 480
rect 48780 400 48832 406
rect 48934 354 49046 480
rect 49988 474 50016 2774
rect 50160 740 50212 746
rect 50160 682 50212 688
rect 50172 480 50200 682
rect 49976 468 50028 474
rect 49976 410 50028 416
rect 48832 348 49046 354
rect 48780 342 49046 348
rect 48792 326 49046 342
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51184 134 51212 2910
rect 52412 2887 52468 2896
rect 51356 2848 51408 2854
rect 53530 2802 53558 3060
rect 54634 2802 54662 3060
rect 55738 2802 55766 3060
rect 56842 2802 56870 3060
rect 57946 2825 57974 3060
rect 51356 2790 51408 2796
rect 51368 480 51396 2790
rect 53484 2774 53558 2802
rect 54588 2774 54662 2802
rect 55692 2774 55766 2802
rect 56796 2774 56870 2802
rect 57932 2816 57988 2825
rect 53010 2680 53066 2689
rect 53010 2615 53066 2624
rect 51172 128 51224 134
rect 51172 70 51224 76
rect 51326 -960 51438 480
rect 52522 354 52634 480
rect 53024 354 53052 2615
rect 53484 1222 53512 2774
rect 53472 1216 53524 1222
rect 53472 1158 53524 1164
rect 52522 326 53052 354
rect 52522 -960 52634 326
rect 53564 128 53616 134
rect 53718 82 53830 480
rect 54588 202 54616 2774
rect 54914 218 55026 480
rect 55692 270 55720 2774
rect 55680 264 55732 270
rect 54914 202 55168 218
rect 55680 206 55732 212
rect 56018 218 56130 480
rect 56796 338 56824 2774
rect 57932 2751 57988 2760
rect 58438 2816 58494 2825
rect 59050 2802 59078 3060
rect 58438 2751 58494 2760
rect 59004 2774 59078 2802
rect 59268 2848 59320 2854
rect 60154 2802 60182 3060
rect 59268 2790 59320 2796
rect 58452 480 58480 2751
rect 59004 1290 59032 2774
rect 59280 1358 59308 2790
rect 60108 2774 60182 2802
rect 60832 2848 60884 2854
rect 61258 2802 61286 3060
rect 62362 2802 62390 3060
rect 63466 2802 63494 3060
rect 60832 2790 60884 2796
rect 59634 2000 59690 2009
rect 59634 1935 59690 1944
rect 59268 1352 59320 1358
rect 59268 1294 59320 1300
rect 58992 1284 59044 1290
rect 58992 1226 59044 1232
rect 59648 480 59676 1935
rect 60108 542 60136 2774
rect 60096 536 60148 542
rect 57214 354 57326 480
rect 57072 338 57326 354
rect 56784 332 56836 338
rect 56784 274 56836 280
rect 57060 332 57326 338
rect 57112 326 57326 332
rect 57060 274 57112 280
rect 56416 264 56468 270
rect 56018 212 56416 218
rect 56018 206 56468 212
rect 54576 196 54628 202
rect 54576 138 54628 144
rect 54914 196 55180 202
rect 54914 190 55128 196
rect 53616 76 53830 82
rect 53564 70 53830 76
rect 53576 54 53830 70
rect 53718 -960 53830 54
rect 54914 -960 55026 190
rect 55128 138 55180 144
rect 56018 190 56456 206
rect 56018 -960 56130 190
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60096 478 60148 484
rect 60844 480 60872 2790
rect 61212 2774 61286 2802
rect 62316 2774 62390 2802
rect 63420 2774 63494 2802
rect 64326 2816 64382 2825
rect 60802 -960 60914 480
rect 61212 105 61240 2774
rect 62316 610 62344 2774
rect 63420 678 63448 2774
rect 64570 2802 64598 3060
rect 64382 2774 64598 2802
rect 65674 2802 65702 3060
rect 66778 2802 66806 3060
rect 67882 2802 67910 3060
rect 68986 2961 69014 3060
rect 68972 2952 69028 2961
rect 68972 2887 69028 2896
rect 65674 2774 65748 2802
rect 64326 2751 64382 2760
rect 65522 2136 65578 2145
rect 65522 2071 65578 2080
rect 63408 672 63460 678
rect 63408 614 63460 620
rect 62304 604 62356 610
rect 62304 546 62356 552
rect 64328 604 64380 610
rect 64328 546 64380 552
rect 63408 536 63460 542
rect 61844 468 61896 474
rect 61844 410 61896 416
rect 61856 354 61884 410
rect 61998 354 62110 480
rect 61856 326 62110 354
rect 61198 96 61254 105
rect 61198 31 61254 40
rect 61998 -960 62110 326
rect 63194 354 63306 480
rect 63408 478 63460 484
rect 64340 480 64368 546
rect 65536 480 65564 2071
rect 63420 354 63448 478
rect 63194 326 63448 354
rect 63194 -960 63306 326
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 65720 406 65748 2774
rect 66732 2774 66806 2802
rect 67836 2774 67910 2802
rect 68928 2848 68980 2854
rect 70090 2802 70118 3060
rect 68928 2790 68980 2796
rect 66732 746 66760 2774
rect 66994 2272 67050 2281
rect 66824 2230 66994 2258
rect 66720 740 66772 746
rect 66720 682 66772 688
rect 66824 626 66852 2230
rect 66994 2207 67050 2216
rect 67836 1358 67864 2774
rect 68940 1358 68968 2790
rect 70044 2774 70118 2802
rect 70308 2848 70360 2854
rect 71194 2802 71222 3060
rect 72298 2802 72326 3060
rect 73402 2802 73430 3060
rect 74506 2961 74534 3060
rect 74492 2952 74548 2961
rect 74492 2887 74548 2896
rect 75610 2802 75638 3060
rect 70308 2790 70360 2796
rect 69110 2408 69166 2417
rect 69110 2343 69166 2352
rect 67824 1352 67876 1358
rect 67824 1294 67876 1300
rect 68928 1352 68980 1358
rect 68928 1294 68980 1300
rect 67916 1216 67968 1222
rect 67916 1158 67968 1164
rect 66732 598 66852 626
rect 66732 480 66760 598
rect 67928 480 67956 1158
rect 69124 480 69152 2343
rect 65708 400 65760 406
rect 65708 342 65760 348
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70044 134 70072 2774
rect 70320 480 70348 2790
rect 71148 2774 71222 2802
rect 72252 2774 72326 2802
rect 73356 2774 73430 2802
rect 75564 2774 75638 2802
rect 76194 2816 76250 2825
rect 70032 128 70084 134
rect 70032 70 70084 76
rect 70278 -960 70390 480
rect 71148 202 71176 2774
rect 71136 196 71188 202
rect 71136 138 71188 144
rect 71474 82 71586 480
rect 72252 270 72280 2774
rect 72606 2544 72662 2553
rect 72606 2479 72662 2488
rect 72620 480 72648 2479
rect 72240 264 72292 270
rect 72240 206 72292 212
rect 71688 128 71740 134
rect 71474 76 71688 82
rect 71474 70 71740 76
rect 71474 54 71728 70
rect 71474 -960 71586 54
rect 72578 -960 72690 480
rect 73356 338 73384 2774
rect 75564 2009 75592 2774
rect 76714 2802 76742 3060
rect 76194 2751 76250 2760
rect 76668 2774 76742 2802
rect 77208 2848 77260 2854
rect 77818 2802 77846 3060
rect 78922 2802 78950 3060
rect 80026 2802 80054 3060
rect 81130 2802 81158 3060
rect 77208 2790 77260 2796
rect 75550 2000 75606 2009
rect 75550 1935 75606 1944
rect 76208 480 76236 2751
rect 76668 1358 76696 2774
rect 76656 1352 76708 1358
rect 76656 1294 76708 1300
rect 77220 1290 77248 2790
rect 77772 2774 77846 2802
rect 78876 2774 78950 2802
rect 79980 2774 80054 2802
rect 81084 2774 81158 2802
rect 82084 2848 82136 2854
rect 82234 2802 82262 3060
rect 83338 2802 83366 3060
rect 84442 2802 84470 3060
rect 85546 2802 85574 3060
rect 86650 2802 86678 3060
rect 87754 2802 87782 3060
rect 88858 2802 88886 3060
rect 89962 2802 89990 3060
rect 91066 2825 91094 3060
rect 82084 2790 82136 2796
rect 77208 1284 77260 1290
rect 77208 1226 77260 1232
rect 77390 640 77446 649
rect 77390 575 77446 584
rect 77404 480 77432 575
rect 73344 332 73396 338
rect 73344 274 73396 280
rect 73774 218 73886 480
rect 73632 202 73886 218
rect 73620 196 73886 202
rect 73672 190 73886 196
rect 73620 138 73672 144
rect 73774 -960 73886 190
rect 74970 218 75082 480
rect 75368 264 75420 270
rect 74970 212 75368 218
rect 74970 206 75420 212
rect 74970 190 75408 206
rect 74970 -960 75082 190
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 77772 474 77800 2774
rect 78876 542 78904 2774
rect 79980 610 80008 2774
rect 81084 2145 81112 2774
rect 81070 2136 81126 2145
rect 81070 2071 81126 2080
rect 81440 1216 81492 1222
rect 81440 1158 81492 1164
rect 79968 604 80020 610
rect 79968 546 80020 552
rect 78864 536 78916 542
rect 77760 468 77812 474
rect 77760 410 77812 416
rect 78404 400 78456 406
rect 78558 354 78670 480
rect 78864 478 78916 484
rect 79662 354 79774 480
rect 78456 348 78670 354
rect 78404 342 78670 348
rect 78416 326 78670 342
rect 79520 338 79774 354
rect 78558 -960 78670 326
rect 79508 332 79774 338
rect 79560 326 79774 332
rect 79508 274 79560 280
rect 79662 -960 79774 326
rect 80858 354 80970 480
rect 81452 354 81480 1158
rect 82096 480 82124 2790
rect 82188 2774 82262 2802
rect 83292 2774 83366 2802
rect 84396 2774 84470 2802
rect 85500 2774 85574 2802
rect 86604 2774 86678 2802
rect 87708 2774 87782 2802
rect 88812 2774 88886 2802
rect 89916 2774 89990 2802
rect 91052 2816 91108 2825
rect 82188 2281 82216 2774
rect 82174 2272 82230 2281
rect 82174 2207 82230 2216
rect 83292 1358 83320 2774
rect 84396 2417 84424 2774
rect 84382 2408 84438 2417
rect 84382 2343 84438 2352
rect 83280 1352 83332 1358
rect 83280 1294 83332 1300
rect 85500 1290 85528 2774
rect 85488 1284 85540 1290
rect 85488 1226 85540 1232
rect 83292 598 83504 626
rect 83292 480 83320 598
rect 83476 513 83504 598
rect 84488 598 84700 626
rect 83462 504 83518 513
rect 80858 326 81480 354
rect 80858 -960 80970 326
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84488 480 84516 598
rect 83462 439 83518 448
rect 84446 -960 84558 480
rect 84672 377 84700 598
rect 84658 368 84714 377
rect 84658 303 84714 312
rect 85642 354 85754 480
rect 86132 468 86184 474
rect 86132 410 86184 416
rect 86144 354 86172 410
rect 85642 326 86172 354
rect 85642 -960 85754 326
rect 86604 134 86632 2774
rect 87708 2553 87736 2774
rect 87694 2544 87750 2553
rect 87694 2479 87750 2488
rect 86592 128 86644 134
rect 86592 70 86644 76
rect 86684 128 86736 134
rect 86838 82 86950 480
rect 87786 368 87842 377
rect 87942 354 88054 480
rect 87842 326 88054 354
rect 87786 303 87842 312
rect 86736 76 86950 82
rect 86684 70 86950 76
rect 86696 54 86950 70
rect 86838 -960 86950 54
rect 87942 -960 88054 326
rect 88812 202 88840 2774
rect 89138 218 89250 480
rect 89916 270 89944 2774
rect 91052 2751 91108 2760
rect 91558 2816 91614 2825
rect 92170 2802 92198 3060
rect 93274 2802 93302 3060
rect 94378 2802 94406 3060
rect 95482 2802 95510 3060
rect 96586 2854 96614 3060
rect 91558 2751 91614 2760
rect 92124 2774 92198 2802
rect 93228 2774 93302 2802
rect 94332 2774 94406 2802
rect 95436 2774 95510 2802
rect 96574 2848 96626 2854
rect 97690 2802 97718 3060
rect 96574 2790 96626 2796
rect 97644 2774 97718 2802
rect 98794 2802 98822 3060
rect 99898 2802 99926 3060
rect 101002 2802 101030 3060
rect 102106 2802 102134 3060
rect 103210 2802 103238 3060
rect 104314 2802 104342 3060
rect 105418 2825 105446 3060
rect 98794 2774 98868 2802
rect 99898 2774 99972 2802
rect 91572 480 91600 2751
rect 92124 649 92152 2774
rect 92110 640 92166 649
rect 92110 575 92166 584
rect 89904 264 89956 270
rect 89138 202 89576 218
rect 89904 206 89956 212
rect 88800 196 88852 202
rect 88800 138 88852 144
rect 89138 196 89588 202
rect 89138 190 89536 196
rect 89138 -960 89250 190
rect 89536 138 89588 144
rect 90178 96 90234 105
rect 90334 82 90446 480
rect 90234 54 90446 82
rect 90178 31 90234 40
rect 90334 -960 90446 54
rect 91530 -960 91642 480
rect 92572 264 92624 270
rect 92726 218 92838 480
rect 93228 406 93256 2774
rect 93950 2000 94006 2009
rect 93950 1935 94006 1944
rect 93964 480 93992 1935
rect 93216 400 93268 406
rect 93216 342 93268 348
rect 92624 212 92838 218
rect 92572 206 92838 212
rect 92584 190 92838 206
rect 92726 -960 92838 190
rect 93922 -960 94034 480
rect 94332 338 94360 2774
rect 95436 1222 95464 2774
rect 95424 1216 95476 1222
rect 95424 1158 95476 1164
rect 97644 513 97672 2774
rect 97908 1216 97960 1222
rect 97908 1158 97960 1164
rect 97630 504 97686 513
rect 95118 354 95230 480
rect 94976 338 95230 354
rect 96068 400 96120 406
rect 96222 354 96334 480
rect 96120 348 96334 354
rect 96068 342 96334 348
rect 94320 332 94372 338
rect 94320 274 94372 280
rect 94964 332 95230 338
rect 95016 326 95230 332
rect 96080 326 96334 342
rect 94964 274 95016 280
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 354 97530 480
rect 97630 439 97686 448
rect 97920 354 97948 1158
rect 98644 672 98696 678
rect 98644 614 98696 620
rect 98656 480 98684 614
rect 98840 513 98868 2774
rect 99746 2272 99802 2281
rect 99746 2207 99802 2216
rect 99760 626 99788 2207
rect 99760 598 99880 626
rect 99944 610 99972 2774
rect 100864 2774 101030 2802
rect 102060 2774 102134 2802
rect 103164 2774 103238 2802
rect 104176 2774 104342 2802
rect 105404 2816 105460 2825
rect 98826 504 98882 513
rect 97418 326 97948 354
rect 97418 -960 97530 326
rect 98614 -960 98726 480
rect 99852 480 99880 598
rect 99932 604 99984 610
rect 99932 546 99984 552
rect 98826 439 98882 448
rect 99810 -960 99922 480
rect 100864 134 100892 2774
rect 101034 2136 101090 2145
rect 101034 2071 101090 2080
rect 101048 480 101076 2071
rect 102060 785 102088 2774
rect 102230 2408 102286 2417
rect 102230 2343 102286 2352
rect 102046 776 102102 785
rect 102046 711 102102 720
rect 102244 480 102272 2343
rect 100852 128 100904 134
rect 100852 70 100904 76
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103164 202 103192 2774
rect 103152 196 103204 202
rect 103152 138 103204 144
rect 103306 82 103418 480
rect 103520 128 103572 134
rect 103306 76 103520 82
rect 104176 105 104204 2774
rect 106522 2802 106550 3060
rect 107626 2802 107654 3060
rect 108730 2802 108758 3060
rect 109834 2802 109862 3060
rect 110938 2802 110966 3060
rect 112042 2802 112070 3060
rect 113146 2802 113174 3060
rect 114250 2802 114278 3060
rect 115354 2802 115382 3060
rect 116458 2802 116486 3060
rect 117562 2802 117590 3060
rect 105404 2751 105460 2760
rect 106476 2774 106550 2802
rect 107580 2774 107654 2802
rect 108684 2774 108758 2802
rect 109788 2774 109862 2802
rect 110892 2774 110966 2802
rect 111996 2774 112070 2802
rect 113100 2774 113174 2802
rect 114204 2774 114278 2802
rect 115308 2774 115382 2802
rect 116228 2774 116486 2802
rect 117516 2774 117590 2802
rect 117686 2816 117742 2825
rect 105726 2544 105782 2553
rect 105726 2479 105782 2488
rect 104532 1352 104584 1358
rect 104532 1294 104584 1300
rect 104544 480 104572 1294
rect 105740 480 105768 2479
rect 103306 70 103572 76
rect 104162 96 104218 105
rect 103306 54 103560 70
rect 103306 -960 103418 54
rect 104162 31 104218 40
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 270 106504 2774
rect 107580 2009 107608 2774
rect 107566 2000 107622 2009
rect 107566 1935 107622 1944
rect 108118 2000 108174 2009
rect 108118 1935 108174 1944
rect 107200 1284 107252 1290
rect 107200 1226 107252 1232
rect 107212 626 107240 1226
rect 106936 598 107240 626
rect 106936 480 106964 598
rect 108132 480 108160 1935
rect 106464 264 106516 270
rect 106464 206 106516 212
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 108684 338 108712 2774
rect 109314 2680 109370 2689
rect 109314 2615 109370 2624
rect 109328 480 109356 2615
rect 108672 332 108724 338
rect 108672 274 108724 280
rect 109286 -960 109398 480
rect 109788 406 109816 2774
rect 110892 1222 110920 2774
rect 111614 1864 111670 1873
rect 111614 1799 111670 1808
rect 110880 1216 110932 1222
rect 110880 1158 110932 1164
rect 110972 1148 111024 1154
rect 110972 1090 111024 1096
rect 109776 400 109828 406
rect 109776 342 109828 348
rect 110482 354 110594 480
rect 110984 354 111012 1090
rect 111628 480 111656 1799
rect 111996 678 112024 2774
rect 113100 2281 113128 2774
rect 113086 2272 113142 2281
rect 113086 2207 113142 2216
rect 114204 2145 114232 2774
rect 115308 2417 115336 2774
rect 115294 2408 115350 2417
rect 115294 2343 115350 2352
rect 114190 2136 114246 2145
rect 114190 2071 114246 2080
rect 115202 2136 115258 2145
rect 115202 2071 115258 2080
rect 112810 1728 112866 1737
rect 112810 1663 112866 1672
rect 111984 672 112036 678
rect 111984 614 112036 620
rect 112824 480 112852 1663
rect 115216 480 115244 2071
rect 110482 326 111012 354
rect 110482 -960 110594 326
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 218 114090 480
rect 113978 202 114416 218
rect 113978 196 114428 202
rect 113978 190 114376 196
rect 113978 -960 114090 190
rect 114376 138 114428 144
rect 115174 -960 115286 480
rect 116228 134 116256 2774
rect 117516 1358 117544 2774
rect 118666 2802 118694 3060
rect 119770 2802 119798 3060
rect 120874 2802 120902 3060
rect 121978 2802 122006 3060
rect 123082 2802 123110 3060
rect 124186 2802 124214 3060
rect 125290 2802 125318 3060
rect 126394 2802 126422 3060
rect 127498 2802 127526 3060
rect 128602 2802 128630 3060
rect 129706 2825 129734 3060
rect 117686 2751 117742 2760
rect 118620 2774 118694 2802
rect 119724 2774 119798 2802
rect 120828 2774 120902 2802
rect 121932 2774 122006 2802
rect 123036 2774 123110 2802
rect 124140 2774 124214 2802
rect 125244 2774 125318 2802
rect 126348 2774 126422 2802
rect 127452 2774 127526 2802
rect 128556 2774 128630 2802
rect 129692 2816 129748 2825
rect 117700 1442 117728 2751
rect 118620 2553 118648 2774
rect 118606 2544 118662 2553
rect 118606 2479 118662 2488
rect 117608 1414 117728 1442
rect 117504 1352 117556 1358
rect 117504 1294 117556 1300
rect 116492 1216 116544 1222
rect 116492 1158 116544 1164
rect 116504 626 116532 1158
rect 116412 598 116532 626
rect 116412 480 116440 598
rect 117608 480 117636 1414
rect 119724 1290 119752 2774
rect 120828 2009 120856 2774
rect 121932 2689 121960 2774
rect 121918 2680 121974 2689
rect 121918 2615 121974 2624
rect 120814 2000 120870 2009
rect 120814 1935 120870 1944
rect 119896 1352 119948 1358
rect 119896 1294 119948 1300
rect 119712 1284 119764 1290
rect 119712 1226 119764 1232
rect 119908 480 119936 1294
rect 121368 1284 121420 1290
rect 121368 1226 121420 1232
rect 121380 626 121408 1226
rect 123036 1154 123064 2774
rect 124140 1873 124168 2774
rect 124126 1864 124182 1873
rect 124126 1799 124182 1808
rect 125244 1737 125272 2774
rect 125230 1728 125286 1737
rect 125230 1663 125286 1672
rect 123024 1148 123076 1154
rect 123024 1090 123076 1096
rect 125140 1148 125192 1154
rect 125140 1090 125192 1096
rect 123482 776 123538 785
rect 123482 711 123538 720
rect 121104 598 121408 626
rect 121104 480 121132 598
rect 123496 480 123524 711
rect 116216 128 116268 134
rect 116216 70 116268 76
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 82 118874 480
rect 119158 96 119214 105
rect 118762 54 119158 82
rect 118762 -960 118874 54
rect 119158 31 119214 40
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 82 122370 480
rect 122564 128 122616 134
rect 122258 76 122564 82
rect 122258 70 122616 76
rect 122258 54 122604 70
rect 122258 -960 122370 54
rect 123454 -960 123566 480
rect 124650 354 124762 480
rect 125152 354 125180 1090
rect 124650 326 125180 354
rect 124650 -960 124762 326
rect 125690 232 125746 241
rect 125846 218 125958 480
rect 125746 190 125958 218
rect 126348 202 126376 2774
rect 127452 2145 127480 2774
rect 127438 2136 127494 2145
rect 127438 2071 127494 2080
rect 128556 1222 128584 2774
rect 130810 2802 130838 3060
rect 131914 2802 131942 3060
rect 133018 2802 133046 3060
rect 134122 2802 134150 3060
rect 134340 2916 134392 2922
rect 134340 2858 134392 2864
rect 129692 2751 129748 2760
rect 130764 2774 130838 2802
rect 131868 2774 131942 2802
rect 132972 2774 133046 2802
rect 133984 2774 134150 2802
rect 128544 1216 128596 1222
rect 128544 1158 128596 1164
rect 129370 912 129426 921
rect 129370 847 129426 856
rect 126992 598 127204 626
rect 126992 480 127020 598
rect 125690 167 125746 176
rect 125846 -960 125958 190
rect 126336 196 126388 202
rect 126336 138 126388 144
rect 126950 -960 127062 480
rect 127176 377 127204 598
rect 129384 480 129412 847
rect 130566 640 130622 649
rect 130566 575 130622 584
rect 130580 480 130608 575
rect 130764 513 130792 2774
rect 131868 1426 131896 2774
rect 131856 1420 131908 1426
rect 131856 1362 131908 1368
rect 132040 1352 132092 1358
rect 132040 1294 132092 1300
rect 132052 762 132080 1294
rect 132972 1290 133000 2774
rect 132960 1284 133012 1290
rect 132960 1226 133012 1232
rect 132774 1048 132830 1057
rect 132774 983 132830 992
rect 131776 734 132080 762
rect 130750 504 130806 513
rect 127162 368 127218 377
rect 127162 303 127218 312
rect 128146 218 128258 480
rect 128146 202 128400 218
rect 128146 196 128412 202
rect 128146 190 128360 196
rect 128146 -960 128258 190
rect 128360 138 128412 144
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131776 480 131804 734
rect 132788 649 132816 983
rect 132774 640 132830 649
rect 132774 575 132830 584
rect 132958 640 133014 649
rect 132958 575 133014 584
rect 132972 480 133000 575
rect 130750 439 130806 448
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 133984 134 134012 2774
rect 134352 1442 134380 2858
rect 135226 2802 135254 3060
rect 136330 2802 136358 3060
rect 137434 2802 137462 3060
rect 138538 2802 138566 3060
rect 139642 2802 139670 3060
rect 140746 2802 140774 3060
rect 141850 2802 141878 3060
rect 142954 2802 142982 3060
rect 144058 2802 144086 3060
rect 145162 2922 145190 3060
rect 145150 2916 145202 2922
rect 145150 2858 145202 2864
rect 146266 2802 146294 3060
rect 134168 1414 134380 1442
rect 135180 2774 135254 2802
rect 136284 2774 136358 2802
rect 137296 2774 137462 2802
rect 138492 2774 138566 2802
rect 139596 2774 139670 2802
rect 140700 2774 140774 2802
rect 141804 2774 141878 2802
rect 142908 2774 142982 2802
rect 144012 2774 144086 2802
rect 146220 2774 146294 2802
rect 147126 2816 147182 2825
rect 134168 480 134196 1414
rect 135180 785 135208 2774
rect 135258 2000 135314 2009
rect 135258 1935 135314 1944
rect 135166 776 135222 785
rect 135166 711 135222 720
rect 135272 480 135300 1935
rect 136284 1222 136312 2774
rect 136272 1216 136324 1222
rect 136272 1158 136324 1164
rect 136454 776 136510 785
rect 136454 711 136510 720
rect 136468 480 136496 711
rect 133972 128 134024 134
rect 133972 70 134024 76
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137296 241 137324 2774
rect 137282 232 137338 241
rect 137282 167 137338 176
rect 137466 232 137522 241
rect 137622 218 137734 480
rect 138492 377 138520 2774
rect 138478 368 138534 377
rect 138478 303 138534 312
rect 137522 190 137734 218
rect 137466 167 137522 176
rect 137622 -960 137734 190
rect 138818 82 138930 480
rect 139596 202 139624 2774
rect 140700 921 140728 2774
rect 141238 2272 141294 2281
rect 141238 2207 141294 2216
rect 140686 912 140742 921
rect 140686 847 140742 856
rect 141252 480 141280 2207
rect 141804 1057 141832 2774
rect 142434 2136 142490 2145
rect 142434 2071 142490 2080
rect 141790 1048 141846 1057
rect 141790 983 141846 992
rect 142448 480 142476 2071
rect 142908 1358 142936 2774
rect 143538 2408 143594 2417
rect 143538 2343 143594 2352
rect 142896 1352 142948 1358
rect 142896 1294 142948 1300
rect 143552 480 143580 2343
rect 144012 649 144040 2774
rect 146220 2009 146248 2774
rect 147370 2802 147398 3060
rect 147126 2751 147182 2760
rect 147324 2774 147398 2802
rect 148474 2802 148502 3060
rect 149578 2802 149606 3060
rect 150682 2802 150710 3060
rect 151786 2802 151814 3060
rect 152890 2802 152918 3060
rect 148474 2774 148548 2802
rect 146206 2000 146262 2009
rect 146206 1935 146262 1944
rect 146208 1352 146260 1358
rect 146208 1294 146260 1300
rect 146220 762 146248 1294
rect 145944 734 146248 762
rect 143998 640 144054 649
rect 143998 575 144054 584
rect 145944 480 145972 734
rect 147140 480 147168 2751
rect 147324 785 147352 2774
rect 148322 2000 148378 2009
rect 148322 1935 148378 1944
rect 147310 776 147366 785
rect 147310 711 147366 720
rect 148336 480 148364 1935
rect 148520 513 148548 2774
rect 149348 2774 149606 2802
rect 150452 2774 150710 2802
rect 151740 2774 151814 2802
rect 152844 2774 152918 2802
rect 153016 2848 153068 2854
rect 153994 2802 154022 3060
rect 155098 2802 155126 3060
rect 156202 2802 156230 3060
rect 157306 2825 157334 3060
rect 153016 2790 153068 2796
rect 148506 504 148562 513
rect 139584 196 139636 202
rect 139584 138 139636 144
rect 139216 128 139268 134
rect 138818 76 139216 82
rect 138818 70 139268 76
rect 139858 96 139914 105
rect 138818 54 139256 70
rect 138818 -960 138930 54
rect 140014 82 140126 480
rect 139914 54 140126 82
rect 139858 31 139914 40
rect 140014 -960 140126 54
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 218 144818 480
rect 144706 202 144960 218
rect 144706 196 144972 202
rect 144706 190 144920 196
rect 144706 -960 144818 190
rect 144920 138 144972 144
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 148506 439 148562 448
rect 149348 134 149376 2774
rect 149518 2544 149574 2553
rect 149518 2479 149574 2488
rect 149532 480 149560 2479
rect 149336 128 149388 134
rect 149336 70 149388 76
rect 149490 -960 149602 480
rect 150346 96 150402 105
rect 150452 82 150480 2774
rect 150622 2680 150678 2689
rect 150622 2615 150678 2624
rect 150636 480 150664 2615
rect 151740 2281 151768 2774
rect 151726 2272 151782 2281
rect 151726 2207 151782 2216
rect 152844 2145 152872 2774
rect 152830 2136 152886 2145
rect 152830 2071 152886 2080
rect 151818 1864 151874 1873
rect 151818 1799 151874 1808
rect 151832 480 151860 1799
rect 153028 480 153056 2790
rect 153948 2774 154022 2802
rect 155052 2774 155126 2802
rect 156156 2774 156230 2802
rect 157292 2816 157348 2825
rect 153948 2417 153976 2774
rect 153934 2408 153990 2417
rect 153934 2343 153990 2352
rect 154210 2136 154266 2145
rect 154210 2071 154266 2080
rect 154224 480 154252 2071
rect 150402 54 150480 82
rect 150346 31 150402 40
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155052 202 155080 2774
rect 155406 2272 155462 2281
rect 155406 2207 155462 2216
rect 155420 480 155448 2207
rect 156156 1358 156184 2774
rect 158410 2802 158438 3060
rect 159514 2802 159542 3060
rect 160618 2802 160646 3060
rect 161722 2802 161750 3060
rect 162826 2854 162854 3060
rect 157292 2751 157348 2760
rect 158364 2774 158438 2802
rect 159468 2774 159542 2802
rect 160572 2774 160646 2802
rect 161676 2774 161750 2802
rect 162814 2848 162866 2854
rect 163930 2802 163958 3060
rect 165034 2802 165062 3060
rect 166138 2802 166166 3060
rect 167242 2802 167270 3060
rect 168346 2802 168374 3060
rect 169450 2802 169478 3060
rect 169576 2916 169628 2922
rect 169576 2858 169628 2864
rect 162814 2790 162866 2796
rect 163884 2774 163958 2802
rect 164988 2774 165062 2802
rect 166092 2774 166166 2802
rect 167196 2774 167270 2802
rect 168024 2774 168374 2802
rect 169404 2774 169478 2802
rect 156602 2408 156658 2417
rect 156602 2343 156658 2352
rect 156144 1352 156196 1358
rect 156144 1294 156196 1300
rect 156616 480 156644 2343
rect 158364 2009 158392 2774
rect 159468 2553 159496 2774
rect 160572 2689 160600 2774
rect 160558 2680 160614 2689
rect 160558 2615 160614 2624
rect 159454 2544 159510 2553
rect 159454 2479 159510 2488
rect 158350 2000 158406 2009
rect 158350 1935 158406 1944
rect 161294 2000 161350 2009
rect 161294 1935 161350 1944
rect 157798 1728 157854 1737
rect 157798 1663 157854 1672
rect 157812 480 157840 1663
rect 160112 598 160324 626
rect 160112 480 160140 598
rect 160296 513 160324 598
rect 160282 504 160338 513
rect 155040 196 155092 202
rect 155040 138 155092 144
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 82 158986 480
rect 159270 96 159326 105
rect 158874 54 159270 82
rect 158874 -960 158986 54
rect 159270 31 159326 40
rect 160070 -960 160182 480
rect 161308 480 161336 1935
rect 161676 1873 161704 2774
rect 162490 2544 162546 2553
rect 162490 2479 162546 2488
rect 161662 1864 161718 1873
rect 161662 1799 161718 1808
rect 162504 480 162532 2479
rect 163884 2145 163912 2774
rect 164988 2281 165016 2774
rect 166092 2417 166120 2774
rect 166078 2408 166134 2417
rect 166078 2343 166134 2352
rect 164974 2272 165030 2281
rect 164974 2207 165030 2216
rect 163870 2136 163926 2145
rect 163870 2071 163926 2080
rect 167196 1737 167224 2774
rect 167182 1728 167238 1737
rect 167182 1663 167238 1672
rect 164148 1352 164200 1358
rect 164148 1294 164200 1300
rect 164882 1320 164938 1329
rect 160282 439 160338 448
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 354 163770 480
rect 164160 354 164188 1294
rect 164882 1255 164938 1264
rect 164896 480 164924 1255
rect 167182 776 167238 785
rect 167182 711 167238 720
rect 165908 598 166120 626
rect 163658 326 164188 354
rect 163658 -960 163770 326
rect 164854 -960 164966 480
rect 165908 377 165936 598
rect 166092 480 166120 598
rect 167196 480 167224 711
rect 165894 368 165950 377
rect 165894 303 165950 312
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168024 105 168052 2774
rect 168378 1048 168434 1057
rect 168378 983 168434 992
rect 168392 480 168420 983
rect 169404 513 169432 2774
rect 169390 504 169446 513
rect 168010 96 168066 105
rect 168010 31 168066 40
rect 168350 -960 168462 480
rect 169588 480 169616 2858
rect 170554 2802 170582 3060
rect 171658 2802 171686 3060
rect 172762 2802 172790 3060
rect 173866 2802 173894 3060
rect 174970 2802 174998 3060
rect 176074 2802 176102 3060
rect 177178 2802 177206 3060
rect 178282 2922 178310 3060
rect 178270 2916 178322 2922
rect 178270 2858 178322 2864
rect 179386 2802 179414 3060
rect 180490 2802 180518 3060
rect 181594 2802 181622 3060
rect 182698 2802 182726 3060
rect 183802 2802 183830 3060
rect 184906 2802 184934 3060
rect 186010 2802 186038 3060
rect 170508 2774 170582 2802
rect 171612 2774 171686 2802
rect 172716 2774 172790 2802
rect 173820 2774 173894 2802
rect 174924 2774 174998 2802
rect 176028 2774 176102 2802
rect 177132 2774 177206 2802
rect 179340 2774 179414 2802
rect 180444 2774 180518 2802
rect 181548 2774 181622 2802
rect 182652 2774 182726 2802
rect 183572 2774 183830 2802
rect 184860 2774 184934 2802
rect 185964 2774 186038 2802
rect 186134 2816 186190 2825
rect 170508 2009 170536 2774
rect 171612 2553 171640 2774
rect 171598 2544 171654 2553
rect 171598 2479 171654 2488
rect 170494 2000 170550 2009
rect 170494 1935 170550 1944
rect 172716 1358 172744 2774
rect 172704 1352 172756 1358
rect 173820 1329 173848 2774
rect 172704 1294 172756 1300
rect 173806 1320 173862 1329
rect 173806 1255 173862 1264
rect 174266 1320 174322 1329
rect 174266 1255 174322 1264
rect 171966 1184 172022 1193
rect 171966 1119 172022 1128
rect 170586 504 170642 513
rect 169390 439 169446 448
rect 169546 -960 169658 480
rect 171980 480 172008 1119
rect 173162 640 173218 649
rect 173162 575 173218 584
rect 173176 480 173204 575
rect 174280 480 174308 1255
rect 170586 439 170642 448
rect 170600 354 170628 439
rect 170742 354 170854 480
rect 170600 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 174924 377 174952 2774
rect 176028 785 176056 2774
rect 177132 1057 177160 2774
rect 177118 1048 177174 1057
rect 177118 983 177174 992
rect 177854 1048 177910 1057
rect 177854 983 177910 992
rect 176014 776 176070 785
rect 176014 711 176070 720
rect 176672 598 176884 626
rect 176672 480 176700 598
rect 174910 368 174966 377
rect 174910 303 174966 312
rect 175434 82 175546 480
rect 175830 96 175886 105
rect 175434 54 175830 82
rect 175434 -960 175546 54
rect 175830 31 175886 40
rect 176630 -960 176742 480
rect 176856 377 176884 598
rect 177868 480 177896 983
rect 179050 776 179106 785
rect 179050 711 179106 720
rect 179064 480 179092 711
rect 179340 513 179368 2774
rect 180246 2000 180302 2009
rect 180246 1935 180302 1944
rect 179326 504 179382 513
rect 176842 368 176898 377
rect 176842 303 176898 312
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180260 480 180288 1935
rect 180444 1193 180472 2774
rect 180430 1184 180486 1193
rect 180430 1119 180486 1128
rect 181442 912 181498 921
rect 181442 847 181498 856
rect 181456 480 181484 847
rect 181548 649 181576 2774
rect 182652 1329 182680 2774
rect 182638 1320 182694 1329
rect 182638 1255 182694 1264
rect 181534 640 181590 649
rect 181534 575 181590 584
rect 179326 439 179382 448
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182362 232 182418 241
rect 182518 218 182630 480
rect 182418 190 182630 218
rect 182362 167 182418 176
rect 182518 -960 182630 190
rect 183466 96 183522 105
rect 183572 82 183600 2774
rect 183742 1184 183798 1193
rect 183742 1119 183798 1128
rect 183756 480 183784 1119
rect 184860 649 184888 2774
rect 184938 1320 184994 1329
rect 184938 1255 184994 1264
rect 184846 640 184902 649
rect 184846 575 184902 584
rect 184952 480 184980 1255
rect 185964 1057 185992 2774
rect 187114 2802 187142 3060
rect 188218 2802 188246 3060
rect 189322 2802 189350 3060
rect 190426 2802 190454 3060
rect 191530 2802 191558 3060
rect 192634 2802 192662 3060
rect 193738 2825 193766 3060
rect 186134 2751 186190 2760
rect 187068 2774 187142 2802
rect 188172 2774 188246 2802
rect 189276 2774 189350 2802
rect 190380 2774 190454 2802
rect 191484 2774 191558 2802
rect 192588 2774 192662 2802
rect 193724 2816 193780 2825
rect 185950 1048 186006 1057
rect 185950 983 186006 992
rect 186148 480 186176 2751
rect 187068 785 187096 2774
rect 188172 2009 188200 2774
rect 188158 2000 188214 2009
rect 188158 1935 188214 1944
rect 189276 921 189304 2774
rect 189722 2000 189778 2009
rect 189722 1935 189778 1944
rect 189262 912 189318 921
rect 189262 847 189318 856
rect 187054 776 187110 785
rect 187054 711 187110 720
rect 189736 480 189764 1935
rect 183522 54 183600 82
rect 183466 31 183522 40
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187146 96 187202 105
rect 187302 82 187414 480
rect 187202 54 187414 82
rect 187146 31 187202 40
rect 187302 -960 187414 54
rect 188498 354 188610 480
rect 188986 368 189042 377
rect 188498 326 188986 354
rect 188498 -960 188610 326
rect 188986 303 189042 312
rect 189694 -960 189806 480
rect 190380 241 190408 2774
rect 191484 1193 191512 2774
rect 192588 1329 192616 2774
rect 194842 2802 194870 3060
rect 195946 2802 195974 3060
rect 197050 2802 197078 3060
rect 198154 2802 198182 3060
rect 199258 2802 199286 3060
rect 200362 2802 200390 3060
rect 201466 2802 201494 3060
rect 202570 2802 202598 3060
rect 203674 2802 203702 3060
rect 204778 2802 204806 3060
rect 205882 2802 205910 3060
rect 206986 2802 207014 3060
rect 208090 2802 208118 3060
rect 209194 2802 209222 3060
rect 210298 2802 210326 3060
rect 211402 2802 211430 3060
rect 212506 2802 212534 3060
rect 213610 2802 213638 3060
rect 214714 2802 214742 3060
rect 215818 2802 215846 3060
rect 193724 2751 193780 2760
rect 194796 2774 194870 2802
rect 195900 2774 195974 2802
rect 197004 2774 197078 2802
rect 198108 2774 198182 2802
rect 199212 2774 199286 2802
rect 200316 2774 200390 2802
rect 201420 2774 201494 2802
rect 202524 2774 202598 2802
rect 203536 2774 203702 2802
rect 204732 2774 204806 2802
rect 205836 2774 205910 2802
rect 206940 2774 207014 2802
rect 208044 2774 208118 2802
rect 209148 2774 209222 2802
rect 210252 2774 210326 2802
rect 211356 2774 211430 2802
rect 212460 2774 212534 2802
rect 213564 2774 213638 2802
rect 214668 2774 214742 2802
rect 215772 2774 215846 2802
rect 216922 2802 216950 3060
rect 218026 2802 218054 3060
rect 219130 2802 219158 3060
rect 220234 2802 220262 3060
rect 221338 2802 221366 3060
rect 222442 2802 222470 3060
rect 223546 2802 223574 3060
rect 224650 2802 224678 3060
rect 225754 2802 225782 3060
rect 226858 2802 226886 3060
rect 227962 2802 227990 3060
rect 229066 2802 229094 3060
rect 230170 2802 230198 3060
rect 231274 2802 231302 3060
rect 232378 2802 232406 3060
rect 233482 2802 233510 3060
rect 234586 2802 234614 3060
rect 235690 2802 235718 3060
rect 236794 2802 236822 3060
rect 237898 2802 237926 3060
rect 239002 2802 239030 3060
rect 240106 2802 240134 3060
rect 241210 2802 241238 3060
rect 242314 2802 242342 3060
rect 243418 2802 243446 3060
rect 244522 2802 244550 3060
rect 245626 2802 245654 3060
rect 246730 2802 246758 3060
rect 247834 2802 247862 3060
rect 248938 2802 248966 3060
rect 250042 2802 250070 3060
rect 251146 2802 251174 3060
rect 252250 2802 252278 3060
rect 253354 2802 253382 3060
rect 254458 2802 254486 3060
rect 255562 2802 255590 3060
rect 256666 2802 256694 3060
rect 257770 2802 257798 3060
rect 258874 2802 258902 3060
rect 259978 2802 260006 3060
rect 261082 2802 261110 3060
rect 262186 2802 262214 3060
rect 263290 2802 263318 3060
rect 264394 2802 264422 3060
rect 265498 2802 265526 3060
rect 266602 2802 266630 3060
rect 267706 2802 267734 3060
rect 268810 2802 268838 3060
rect 269914 2802 269942 3060
rect 271018 2802 271046 3060
rect 272122 2802 272150 3060
rect 273226 2802 273254 3060
rect 274330 2802 274358 3060
rect 275434 2802 275462 3060
rect 276538 2802 276566 3060
rect 277642 2802 277670 3060
rect 278746 2802 278774 3060
rect 279850 2802 279878 3060
rect 280954 2802 280982 3060
rect 282058 2802 282086 3060
rect 283162 2938 283190 3060
rect 284266 2938 284294 3060
rect 283162 2910 283236 2938
rect 216922 2774 216996 2802
rect 192574 1320 192630 1329
rect 192574 1255 192630 1264
rect 191470 1184 191526 1193
rect 191470 1119 191526 1128
rect 194414 1184 194470 1193
rect 194414 1119 194470 1128
rect 193218 1048 193274 1057
rect 193218 983 193274 992
rect 192022 912 192078 921
rect 192022 847 192078 856
rect 190826 776 190882 785
rect 190826 711 190882 720
rect 190840 480 190868 711
rect 192036 480 192064 847
rect 193232 480 193260 983
rect 194428 480 194456 1119
rect 190366 232 190422 241
rect 190366 167 190422 176
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 194796 105 194824 2774
rect 195610 1320 195666 1329
rect 195610 1255 195666 1264
rect 195624 480 195652 1255
rect 195900 649 195928 2774
rect 197004 2009 197032 2774
rect 196990 2000 197046 2009
rect 196990 1935 197046 1944
rect 198108 785 198136 2774
rect 199212 921 199240 2774
rect 200316 1057 200344 2774
rect 200486 1728 200542 1737
rect 200408 1686 200486 1714
rect 200302 1048 200358 1057
rect 200302 983 200358 992
rect 199198 912 199254 921
rect 200408 898 200436 1686
rect 200486 1663 200542 1672
rect 201420 1193 201448 2774
rect 201498 1456 201554 1465
rect 201498 1391 201554 1400
rect 201406 1184 201462 1193
rect 201406 1119 201462 1128
rect 199198 847 199254 856
rect 200316 870 200436 898
rect 198094 776 198150 785
rect 198094 711 198150 720
rect 199106 776 199162 785
rect 199106 711 199162 720
rect 195886 640 195942 649
rect 195886 575 195942 584
rect 199120 480 199148 711
rect 200316 480 200344 870
rect 201512 480 201540 1391
rect 202524 1329 202552 2774
rect 202510 1320 202566 1329
rect 202510 1255 202566 1264
rect 202694 1048 202750 1057
rect 202694 983 202750 992
rect 202708 480 202736 983
rect 194782 96 194838 105
rect 194782 31 194838 40
rect 195582 -960 195694 480
rect 196778 82 196890 480
rect 197882 354 197994 480
rect 198370 368 198426 377
rect 197882 326 198370 354
rect 197174 96 197230 105
rect 196778 54 197174 82
rect 196778 -960 196890 54
rect 197174 31 197230 40
rect 197882 -960 197994 326
rect 198370 303 198426 312
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203536 105 203564 2774
rect 203890 1184 203946 1193
rect 203890 1119 203946 1128
rect 203904 480 203932 1119
rect 203522 96 203578 105
rect 203522 31 203578 40
rect 203862 -960 203974 480
rect 204732 377 204760 2774
rect 205086 1320 205142 1329
rect 205086 1255 205142 1264
rect 205100 480 205128 1255
rect 205836 785 205864 2774
rect 206940 1737 206968 2774
rect 207386 2136 207442 2145
rect 207386 2071 207442 2080
rect 206926 1728 206982 1737
rect 206926 1663 206982 1672
rect 206190 1592 206246 1601
rect 206190 1527 206246 1536
rect 205822 776 205878 785
rect 205822 711 205878 720
rect 206204 480 206232 1527
rect 207400 480 207428 2071
rect 208044 1465 208072 2774
rect 208582 2000 208638 2009
rect 208582 1935 208638 1944
rect 208030 1456 208086 1465
rect 208030 1391 208086 1400
rect 208596 480 208624 1935
rect 209148 1057 209176 2774
rect 209778 2272 209834 2281
rect 209778 2207 209834 2216
rect 209134 1048 209190 1057
rect 209134 983 209190 992
rect 209792 480 209820 2207
rect 210252 1193 210280 2774
rect 211356 1329 211384 2774
rect 212170 1864 212226 1873
rect 212170 1799 212226 1808
rect 211342 1320 211398 1329
rect 211342 1255 211398 1264
rect 210238 1184 210294 1193
rect 210238 1119 210294 1128
rect 210974 1184 211030 1193
rect 210974 1119 211030 1128
rect 210988 480 211016 1119
rect 212184 480 212212 1799
rect 212460 1601 212488 2774
rect 213564 2145 213592 2774
rect 213550 2136 213606 2145
rect 213550 2071 213606 2080
rect 214668 2009 214696 2774
rect 215772 2281 215800 2774
rect 216862 2408 216918 2417
rect 216862 2343 216918 2352
rect 215758 2272 215814 2281
rect 215758 2207 215814 2216
rect 214654 2000 214710 2009
rect 214654 1935 214710 1944
rect 213366 1728 213422 1737
rect 213366 1663 213422 1672
rect 212446 1592 212502 1601
rect 212446 1527 212502 1536
rect 213380 480 213408 1663
rect 215666 1592 215722 1601
rect 215666 1527 215722 1536
rect 214470 1456 214526 1465
rect 214470 1391 214526 1400
rect 214484 480 214512 1391
rect 215680 480 215708 1527
rect 216876 480 216904 2343
rect 216968 1193 216996 2774
rect 217980 2774 218054 2802
rect 219084 2774 219158 2802
rect 220188 2774 220262 2802
rect 221292 2774 221366 2802
rect 222396 2774 222470 2802
rect 223500 2774 223574 2802
rect 224604 2774 224678 2802
rect 225708 2774 225782 2802
rect 226812 2774 226886 2802
rect 227916 2774 227990 2802
rect 229020 2774 229094 2802
rect 230124 2774 230198 2802
rect 231228 2774 231302 2802
rect 232332 2774 232406 2802
rect 233436 2774 233510 2802
rect 234540 2774 234614 2802
rect 235644 2774 235718 2802
rect 236748 2774 236822 2802
rect 237852 2774 237926 2802
rect 238956 2774 239030 2802
rect 240060 2774 240134 2802
rect 241164 2774 241238 2802
rect 242268 2774 242342 2802
rect 243372 2774 243446 2802
rect 244476 2774 244550 2802
rect 245580 2774 245654 2802
rect 246684 2774 246758 2802
rect 247788 2774 247862 2802
rect 248892 2774 248966 2802
rect 249996 2774 250070 2802
rect 251100 2774 251174 2802
rect 252204 2774 252278 2802
rect 253308 2774 253382 2802
rect 254412 2774 254486 2802
rect 255516 2774 255590 2802
rect 256620 2774 256694 2802
rect 257724 2774 257798 2802
rect 258828 2774 258902 2802
rect 259932 2774 260006 2802
rect 261036 2774 261110 2802
rect 262140 2774 262214 2802
rect 263244 2774 263318 2802
rect 264348 2774 264422 2802
rect 265452 2774 265526 2802
rect 266556 2774 266630 2802
rect 267660 2774 267734 2802
rect 268764 2774 268838 2802
rect 269868 2774 269942 2802
rect 270972 2774 271046 2802
rect 272076 2774 272150 2802
rect 273180 2774 273254 2802
rect 274284 2774 274358 2802
rect 275388 2774 275462 2802
rect 276492 2774 276566 2802
rect 277596 2774 277670 2802
rect 278700 2774 278774 2802
rect 279804 2774 279878 2802
rect 280908 2774 280982 2802
rect 282012 2774 282086 2802
rect 217980 1873 218008 2774
rect 218058 2680 218114 2689
rect 218058 2615 218114 2624
rect 217966 1864 218022 1873
rect 217966 1799 218022 1808
rect 216954 1184 217010 1193
rect 216954 1119 217010 1128
rect 218072 480 218100 2615
rect 219084 1737 219112 2774
rect 219254 2272 219310 2281
rect 219254 2207 219310 2216
rect 219070 1728 219126 1737
rect 219070 1663 219126 1672
rect 219268 480 219296 2207
rect 220188 1465 220216 2774
rect 220450 2000 220506 2009
rect 220450 1935 220506 1944
rect 220174 1456 220230 1465
rect 220174 1391 220230 1400
rect 220464 480 220492 1935
rect 221292 1601 221320 2774
rect 222396 2417 222424 2774
rect 223500 2689 223528 2774
rect 223486 2680 223542 2689
rect 223486 2615 223542 2624
rect 222382 2408 222438 2417
rect 222382 2343 222438 2352
rect 224604 2281 224632 2774
rect 224590 2272 224646 2281
rect 224590 2207 224646 2216
rect 223946 2136 224002 2145
rect 223946 2071 224002 2080
rect 221554 1864 221610 1873
rect 221554 1799 221610 1808
rect 221278 1592 221334 1601
rect 221278 1527 221334 1536
rect 221568 480 221596 1799
rect 222750 1728 222806 1737
rect 222750 1663 222806 1672
rect 222764 480 222792 1663
rect 223960 480 223988 2071
rect 225708 2009 225736 2774
rect 225694 2000 225750 2009
rect 225694 1935 225750 1944
rect 226812 1873 226840 2774
rect 227534 2000 227590 2009
rect 227534 1935 227590 1944
rect 226798 1864 226854 1873
rect 226798 1799 226854 1808
rect 226338 1592 226394 1601
rect 226338 1527 226394 1536
rect 225142 1456 225198 1465
rect 225142 1391 225198 1400
rect 225156 480 225184 1391
rect 226352 480 226380 1527
rect 227548 480 227576 1935
rect 227916 1737 227944 2774
rect 228730 2408 228786 2417
rect 228730 2343 228786 2352
rect 227902 1728 227958 1737
rect 227902 1663 227958 1672
rect 228744 480 228772 2343
rect 229020 2145 229048 2774
rect 229006 2136 229062 2145
rect 229006 2071 229062 2080
rect 229834 2136 229890 2145
rect 229834 2071 229890 2080
rect 229848 480 229876 2071
rect 230124 1465 230152 2774
rect 231228 1601 231256 2774
rect 232332 2009 232360 2774
rect 233436 2417 233464 2774
rect 233422 2408 233478 2417
rect 233422 2343 233478 2352
rect 234540 2145 234568 2774
rect 234526 2136 234582 2145
rect 234526 2071 234582 2080
rect 232318 2000 232374 2009
rect 232318 1935 232374 1944
rect 233422 1864 233478 1873
rect 233422 1799 233478 1808
rect 231214 1592 231270 1601
rect 231214 1527 231270 1536
rect 232226 1592 232282 1601
rect 232226 1527 232282 1536
rect 230110 1456 230166 1465
rect 230110 1391 230166 1400
rect 231030 1456 231086 1465
rect 231030 1391 231086 1400
rect 231044 480 231072 1391
rect 232240 480 232268 1527
rect 233436 480 233464 1799
rect 234618 1728 234674 1737
rect 234618 1663 234674 1672
rect 234632 480 234660 1663
rect 235644 1465 235672 2774
rect 236748 1601 236776 2774
rect 237852 1873 237880 2774
rect 238114 2000 238170 2009
rect 238114 1935 238170 1944
rect 237838 1864 237894 1873
rect 237838 1799 237894 1808
rect 236734 1592 236790 1601
rect 236734 1527 236790 1536
rect 237010 1592 237066 1601
rect 237010 1527 237066 1536
rect 235630 1456 235686 1465
rect 235630 1391 235686 1400
rect 235814 1456 235870 1465
rect 235814 1391 235870 1400
rect 235828 480 235856 1391
rect 237024 480 237052 1527
rect 238128 480 238156 1935
rect 238956 1737 238984 2774
rect 239310 2136 239366 2145
rect 239310 2071 239366 2080
rect 238942 1728 238998 1737
rect 238942 1663 238998 1672
rect 239324 480 239352 2071
rect 240060 1465 240088 2774
rect 241164 1601 241192 2774
rect 242268 2009 242296 2774
rect 243372 2145 243400 2774
rect 243358 2136 243414 2145
rect 243358 2071 243414 2080
rect 242254 2000 242310 2009
rect 242254 1935 242310 1944
rect 241702 1864 241758 1873
rect 241702 1799 241758 1808
rect 241150 1592 241206 1601
rect 241150 1527 241206 1536
rect 240046 1456 240102 1465
rect 240046 1391 240102 1400
rect 240506 1456 240562 1465
rect 240506 1391 240562 1400
rect 240520 480 240548 1391
rect 241716 480 241744 1799
rect 242898 1728 242954 1737
rect 242898 1663 242954 1672
rect 242912 480 242940 1663
rect 244094 1592 244150 1601
rect 244094 1527 244150 1536
rect 244108 480 244136 1527
rect 244476 1465 244504 2774
rect 245580 1873 245608 2774
rect 246394 2408 246450 2417
rect 246394 2343 246450 2352
rect 245566 1864 245622 1873
rect 245566 1799 245622 1808
rect 244462 1456 244518 1465
rect 244462 1391 244518 1400
rect 245198 1456 245254 1465
rect 245198 1391 245254 1400
rect 245212 480 245240 1391
rect 246408 480 246436 2343
rect 246684 1737 246712 2774
rect 247590 1864 247646 1873
rect 247590 1799 247646 1808
rect 246670 1728 246726 1737
rect 246670 1663 246726 1672
rect 247604 480 247632 1799
rect 247788 1601 247816 2774
rect 248786 2000 248842 2009
rect 248786 1935 248842 1944
rect 247774 1592 247830 1601
rect 247774 1527 247830 1536
rect 248800 480 248828 1935
rect 248892 1465 248920 2774
rect 249996 2417 250024 2774
rect 249982 2408 250038 2417
rect 249982 2343 250038 2352
rect 251100 1873 251128 2774
rect 252204 2009 252232 2774
rect 252190 2000 252246 2009
rect 252190 1935 252246 1944
rect 251086 1864 251142 1873
rect 251086 1799 251142 1808
rect 251178 1728 251234 1737
rect 251178 1663 251234 1672
rect 249982 1592 250038 1601
rect 249982 1527 250038 1536
rect 248878 1456 248934 1465
rect 248878 1391 248934 1400
rect 249996 480 250024 1527
rect 251192 480 251220 1663
rect 253308 1601 253336 2774
rect 254412 1737 254440 2774
rect 254398 1728 254454 1737
rect 254398 1663 254454 1672
rect 254674 1728 254730 1737
rect 254674 1663 254730 1672
rect 253294 1592 253350 1601
rect 253294 1527 253350 1536
rect 253478 1592 253534 1601
rect 253478 1527 253534 1536
rect 252374 1456 252430 1465
rect 252374 1391 252430 1400
rect 252388 480 252416 1391
rect 253492 480 253520 1527
rect 254688 480 254716 1663
rect 255516 1465 255544 2774
rect 256620 1601 256648 2774
rect 257724 1737 257752 2774
rect 257710 1728 257766 1737
rect 257710 1663 257766 1672
rect 258262 1728 258318 1737
rect 258262 1663 258318 1672
rect 256606 1592 256662 1601
rect 256606 1527 256662 1536
rect 257066 1592 257122 1601
rect 257066 1527 257122 1536
rect 255502 1456 255558 1465
rect 255502 1391 255558 1400
rect 255870 1456 255926 1465
rect 255870 1391 255926 1400
rect 255884 480 255912 1391
rect 257080 480 257108 1527
rect 258276 480 258304 1663
rect 258828 1465 258856 2774
rect 259932 1601 259960 2774
rect 261036 1737 261064 2774
rect 261022 1728 261078 1737
rect 261022 1663 261078 1672
rect 261758 1728 261814 1737
rect 261758 1663 261814 1672
rect 259918 1592 259974 1601
rect 259918 1527 259974 1536
rect 260654 1592 260710 1601
rect 260654 1527 260710 1536
rect 258814 1456 258870 1465
rect 258814 1391 258870 1400
rect 259458 1320 259514 1329
rect 259458 1255 259514 1264
rect 259472 480 259500 1255
rect 260668 480 260696 1527
rect 261772 480 261800 1663
rect 262140 1329 262168 2774
rect 263244 1601 263272 2774
rect 264348 1737 264376 2774
rect 264334 1728 264390 1737
rect 264334 1663 264390 1672
rect 263230 1592 263286 1601
rect 263230 1527 263286 1536
rect 264150 1592 264206 1601
rect 264150 1527 264206 1536
rect 262954 1456 263010 1465
rect 262954 1391 263010 1400
rect 262126 1320 262182 1329
rect 262126 1255 262182 1264
rect 262968 480 262996 1391
rect 264164 480 264192 1527
rect 265452 1465 265480 2774
rect 266556 1601 266584 2774
rect 266542 1592 266598 1601
rect 266542 1527 266598 1536
rect 265438 1456 265494 1465
rect 265438 1391 265494 1400
rect 266542 1184 266598 1193
rect 266542 1119 266598 1128
rect 265346 1048 265402 1057
rect 265346 983 265402 992
rect 265360 480 265388 983
rect 266556 480 266584 1119
rect 267660 1057 267688 2774
rect 267738 1320 267794 1329
rect 267738 1255 267794 1264
rect 267646 1048 267702 1057
rect 267646 983 267702 992
rect 267752 480 267780 1255
rect 268764 1193 268792 2774
rect 268842 1456 268898 1465
rect 268842 1391 268898 1400
rect 268750 1184 268806 1193
rect 268750 1119 268806 1128
rect 268856 480 268884 1391
rect 269868 1329 269896 2774
rect 270038 1592 270094 1601
rect 270038 1527 270094 1536
rect 269854 1320 269910 1329
rect 269854 1255 269910 1264
rect 270052 480 270080 1527
rect 270972 1465 271000 2774
rect 272076 1601 272104 2774
rect 272062 1592 272118 1601
rect 272062 1527 272118 1536
rect 270958 1456 271014 1465
rect 270958 1391 271014 1400
rect 273180 1329 273208 2774
rect 271234 1320 271290 1329
rect 271234 1255 271290 1264
rect 273166 1320 273222 1329
rect 273166 1255 273222 1264
rect 273626 1320 273682 1329
rect 273626 1255 273682 1264
rect 271248 480 271276 1255
rect 272430 1184 272486 1193
rect 272430 1119 272486 1128
rect 272444 480 272472 1119
rect 273640 480 273668 1255
rect 274284 1193 274312 2774
rect 275388 1329 275416 2774
rect 275374 1320 275430 1329
rect 275374 1255 275430 1264
rect 276018 1320 276074 1329
rect 276018 1255 276074 1264
rect 274270 1184 274326 1193
rect 274270 1119 274326 1128
rect 274822 1184 274878 1193
rect 274822 1119 274878 1128
rect 274836 480 274864 1119
rect 276032 480 276060 1255
rect 276492 1193 276520 2774
rect 277596 1329 277624 2774
rect 277582 1320 277638 1329
rect 277582 1255 277638 1264
rect 278700 1193 278728 2774
rect 279514 1320 279570 1329
rect 279514 1255 279570 1264
rect 276478 1184 276534 1193
rect 276478 1119 276534 1128
rect 277122 1184 277178 1193
rect 277122 1119 277178 1128
rect 278686 1184 278742 1193
rect 278686 1119 278742 1128
rect 277136 480 277164 1119
rect 278318 1048 278374 1057
rect 278318 983 278374 992
rect 278332 480 278360 983
rect 279528 480 279556 1255
rect 279804 1057 279832 2774
rect 280908 1329 280936 2774
rect 280894 1320 280950 1329
rect 280894 1255 280950 1264
rect 281906 1320 281962 1329
rect 281906 1255 281962 1264
rect 280710 1184 280766 1193
rect 280710 1119 280766 1128
rect 279790 1048 279846 1057
rect 279790 983 279846 992
rect 280724 480 280752 1119
rect 281920 480 281948 1255
rect 282012 1193 282040 2774
rect 283208 1329 283236 2910
rect 283300 2910 284294 2938
rect 283194 1320 283250 1329
rect 283194 1255 283250 1264
rect 281998 1184 282054 1193
rect 283300 1170 283328 2910
rect 285370 2802 285398 3060
rect 286474 2802 286502 3060
rect 287578 2802 287606 3060
rect 288682 2802 288710 3060
rect 289786 2802 289814 3060
rect 290890 2802 290918 3060
rect 291994 2802 292022 3060
rect 293098 2802 293126 3060
rect 294202 2802 294230 3060
rect 295306 2802 295334 3060
rect 296410 2802 296438 3060
rect 297514 2802 297542 3060
rect 298618 2802 298646 3060
rect 299722 2802 299750 3060
rect 300826 2802 300854 3060
rect 281998 1119 282054 1128
rect 283116 1142 283328 1170
rect 284312 2774 285398 2802
rect 286428 2774 286502 2802
rect 287532 2774 287606 2802
rect 288636 2774 288710 2802
rect 289464 2774 289814 2802
rect 290200 2774 290918 2802
rect 291856 2774 292022 2802
rect 292592 2774 293126 2802
rect 293696 2774 294230 2802
rect 295260 2774 295334 2802
rect 296088 2774 296438 2802
rect 297468 2774 297542 2802
rect 298480 2774 298646 2802
rect 299676 2774 299750 2802
rect 300780 2774 300854 2802
rect 301930 2802 301958 3060
rect 303034 2802 303062 3060
rect 304138 2802 304166 3060
rect 305242 2802 305270 3060
rect 306346 2802 306374 3060
rect 307450 2802 307478 3060
rect 308554 2802 308582 3060
rect 309658 2802 309686 3060
rect 310762 2802 310790 3060
rect 311866 2802 311894 3060
rect 312970 2802 312998 3060
rect 314074 2802 314102 3060
rect 315178 2802 315206 3060
rect 316282 2802 316310 3060
rect 317386 2938 317414 3060
rect 317386 2910 317460 2938
rect 301930 2774 302004 2802
rect 303034 2774 303200 2802
rect 304138 2774 304212 2802
rect 305242 2774 305592 2802
rect 306346 2774 306420 2802
rect 307450 2774 307984 2802
rect 308554 2774 309088 2802
rect 309658 2774 309824 2802
rect 310762 2774 311480 2802
rect 311866 2774 312216 2802
rect 312970 2774 313044 2802
rect 314074 2774 314148 2802
rect 315178 2774 315252 2802
rect 316282 2774 317368 2802
rect 283116 480 283144 1142
rect 284312 480 284340 2774
rect 286428 1329 286456 2774
rect 287532 1329 287560 2774
rect 288636 1329 288664 2774
rect 285402 1320 285458 1329
rect 285402 1255 285458 1264
rect 286414 1320 286470 1329
rect 286414 1255 286470 1264
rect 286598 1320 286654 1329
rect 286598 1255 286654 1264
rect 287518 1320 287574 1329
rect 287518 1255 287574 1264
rect 287794 1320 287850 1329
rect 287794 1255 287850 1264
rect 288622 1320 288678 1329
rect 288622 1255 288678 1264
rect 285416 480 285444 1255
rect 286612 480 286640 1255
rect 287808 480 287836 1255
rect 204718 368 204774 377
rect 204718 303 204774 312
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 354 289074 480
rect 289464 354 289492 2774
rect 290200 480 290228 2774
rect 288962 326 289492 354
rect 288962 -960 289074 326
rect 290158 -960 290270 480
rect 291354 354 291466 480
rect 291856 354 291884 2774
rect 292592 480 292620 2774
rect 293696 480 293724 2774
rect 291354 326 291884 354
rect 291354 -960 291466 326
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 354 294962 480
rect 295260 354 295288 2774
rect 296088 480 296116 2774
rect 294850 326 295288 354
rect 294850 -960 294962 326
rect 296046 -960 296158 480
rect 297242 354 297354 480
rect 297468 354 297496 2774
rect 298480 480 298508 2774
rect 299676 480 299704 2774
rect 300780 480 300808 2774
rect 301976 480 302004 2774
rect 303172 480 303200 2774
rect 297242 326 297496 354
rect 297242 -960 297354 326
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304184 354 304212 2774
rect 305564 480 305592 2774
rect 304326 354 304438 480
rect 304184 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 2774
rect 307956 480 307984 2774
rect 309060 480 309088 2774
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 2774
rect 311452 480 311480 2774
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 2774
rect 313016 1329 313044 2774
rect 314120 1329 314148 2774
rect 315224 1329 315252 2774
rect 313002 1320 313058 1329
rect 313002 1255 313058 1264
rect 313830 1320 313886 1329
rect 313830 1255 313886 1264
rect 314106 1320 314162 1329
rect 314106 1255 314162 1264
rect 315026 1320 315082 1329
rect 315026 1255 315082 1264
rect 315210 1320 315266 1329
rect 315210 1255 315266 1264
rect 316222 1320 316278 1329
rect 316222 1255 316278 1264
rect 313844 480 313872 1255
rect 315040 480 315068 1255
rect 316236 480 316264 1255
rect 317340 480 317368 2774
rect 317432 1329 317460 2910
rect 318490 2802 318518 3060
rect 318444 2774 318518 2802
rect 319594 2802 319622 3060
rect 320698 2802 320726 3060
rect 321802 2802 321830 3060
rect 322906 2802 322934 3060
rect 319594 2774 319668 2802
rect 320698 2774 320772 2802
rect 321802 2774 321876 2802
rect 317418 1320 317474 1329
rect 317418 1255 317474 1264
rect 318444 1193 318472 2774
rect 319640 1329 319668 2774
rect 318522 1320 318578 1329
rect 318522 1255 318578 1264
rect 319626 1320 319682 1329
rect 319626 1255 319682 1264
rect 318430 1184 318486 1193
rect 318430 1119 318486 1128
rect 318536 480 318564 1255
rect 320744 1193 320772 2774
rect 320914 1320 320970 1329
rect 320914 1255 320970 1264
rect 319718 1184 319774 1193
rect 319718 1119 319774 1128
rect 320730 1184 320786 1193
rect 320730 1119 320786 1128
rect 319732 480 319760 1119
rect 320928 480 320956 1255
rect 321848 1057 321876 2774
rect 322860 2774 322934 2802
rect 324010 2802 324038 3060
rect 325114 2802 325142 3060
rect 326218 2802 326246 3060
rect 327322 2802 327350 3060
rect 328426 2802 328454 3060
rect 324010 2774 324084 2802
rect 325114 2774 325188 2802
rect 326218 2774 326292 2802
rect 327322 2774 327396 2802
rect 322860 1329 322888 2774
rect 322846 1320 322902 1329
rect 322846 1255 322902 1264
rect 324056 1193 324084 2774
rect 325160 1329 325188 2774
rect 324410 1320 324466 1329
rect 324410 1255 324466 1264
rect 325146 1320 325202 1329
rect 325146 1255 325202 1264
rect 322110 1184 322166 1193
rect 322110 1119 322166 1128
rect 324042 1184 324098 1193
rect 324042 1119 324098 1128
rect 321834 1048 321890 1057
rect 321834 983 321890 992
rect 322124 480 322152 1119
rect 323306 1048 323362 1057
rect 323306 983 323362 992
rect 323320 480 323348 983
rect 324424 480 324452 1255
rect 326264 1193 326292 2774
rect 327368 1329 327396 2774
rect 328380 2774 328454 2802
rect 329530 2802 329558 3060
rect 330634 2802 330662 3060
rect 331738 2802 331766 3060
rect 332842 2802 332870 3060
rect 333946 2802 333974 3060
rect 329530 2774 329604 2802
rect 330634 2774 330708 2802
rect 331738 2774 331812 2802
rect 332842 2774 332916 2802
rect 326802 1320 326858 1329
rect 326802 1255 326858 1264
rect 327354 1320 327410 1329
rect 327354 1255 327410 1264
rect 325606 1184 325662 1193
rect 325606 1119 325662 1128
rect 326250 1184 326306 1193
rect 326250 1119 326306 1128
rect 325620 480 325648 1119
rect 326816 480 326844 1255
rect 328380 1193 328408 2774
rect 329576 1329 329604 2774
rect 329194 1320 329250 1329
rect 329194 1255 329250 1264
rect 329562 1320 329618 1329
rect 329562 1255 329618 1264
rect 327998 1184 328054 1193
rect 327998 1119 328054 1128
rect 328366 1184 328422 1193
rect 328366 1119 328422 1128
rect 328012 480 328040 1119
rect 329208 480 329236 1255
rect 330680 1193 330708 2774
rect 331586 1320 331642 1329
rect 331586 1255 331642 1264
rect 330390 1184 330446 1193
rect 330390 1119 330446 1128
rect 330666 1184 330722 1193
rect 330666 1119 330722 1128
rect 330404 480 330432 1119
rect 331600 480 331628 1255
rect 331784 921 331812 2774
rect 332888 1193 332916 2774
rect 333900 2774 333974 2802
rect 335050 2802 335078 3060
rect 336154 2802 336182 3060
rect 337258 2802 337286 3060
rect 338362 2802 338390 3060
rect 339466 2802 339494 3060
rect 335050 2774 335124 2802
rect 336154 2774 336228 2802
rect 337258 2774 337332 2802
rect 338362 2774 338436 2802
rect 332690 1184 332746 1193
rect 332690 1119 332746 1128
rect 332874 1184 332930 1193
rect 332874 1119 332930 1128
rect 331770 912 331826 921
rect 331770 847 331826 856
rect 332704 480 332732 1119
rect 333900 1057 333928 2774
rect 335096 1329 335124 2774
rect 335082 1320 335138 1329
rect 335082 1255 335138 1264
rect 336200 1193 336228 2774
rect 335082 1184 335138 1193
rect 335082 1119 335138 1128
rect 336186 1184 336242 1193
rect 336186 1119 336242 1128
rect 333886 1048 333942 1057
rect 333886 983 333942 992
rect 333886 912 333942 921
rect 333886 847 333942 856
rect 333900 480 333928 847
rect 335096 480 335124 1119
rect 337304 1057 337332 2774
rect 338408 1329 338436 2774
rect 339420 2774 339494 2802
rect 340570 2802 340598 3060
rect 341674 2802 341702 3060
rect 342778 2802 342806 3060
rect 343882 2802 343910 3060
rect 344986 2825 345014 3060
rect 346090 2825 346118 3060
rect 344972 2816 345028 2825
rect 340570 2774 340644 2802
rect 341674 2774 341748 2802
rect 342778 2774 342852 2802
rect 343882 2774 343956 2802
rect 337474 1320 337530 1329
rect 337474 1255 337530 1264
rect 338394 1320 338450 1329
rect 338394 1255 338450 1264
rect 336278 1048 336334 1057
rect 336278 983 336334 992
rect 337290 1048 337346 1057
rect 337290 983 337346 992
rect 336292 480 336320 983
rect 337488 480 337516 1255
rect 339420 1193 339448 2774
rect 338670 1184 338726 1193
rect 338670 1119 338726 1128
rect 339406 1184 339462 1193
rect 339406 1119 339462 1128
rect 338684 480 338712 1119
rect 340616 1057 340644 2774
rect 341720 1329 341748 2774
rect 340970 1320 341026 1329
rect 340970 1255 341026 1264
rect 341706 1320 341762 1329
rect 341706 1255 341762 1264
rect 339866 1048 339922 1057
rect 339866 983 339922 992
rect 340602 1048 340658 1057
rect 340602 983 340658 992
rect 339880 480 339908 983
rect 340984 480 341012 1255
rect 342824 1193 342852 2774
rect 342166 1184 342222 1193
rect 342166 1119 342222 1128
rect 342810 1184 342866 1193
rect 342810 1119 342866 1128
rect 342180 480 342208 1119
rect 343928 1057 343956 2774
rect 344972 2751 345028 2760
rect 346076 2816 346132 2825
rect 347194 2802 347222 3060
rect 348298 2802 348326 3060
rect 349250 2816 349306 2825
rect 347194 2774 347268 2802
rect 348298 2774 348372 2802
rect 346076 2751 346132 2760
rect 347240 1329 347268 2774
rect 347778 2680 347834 2689
rect 347834 2638 348096 2666
rect 347778 2615 347834 2624
rect 344558 1320 344614 1329
rect 344558 1255 344614 1264
rect 347226 1320 347282 1329
rect 347226 1255 347282 1264
rect 343362 1048 343418 1057
rect 343362 983 343418 992
rect 343914 1048 343970 1057
rect 343914 983 343970 992
rect 343376 480 343404 983
rect 344572 480 344600 1255
rect 345754 1184 345810 1193
rect 345754 1119 345810 1128
rect 345768 480 345796 1119
rect 346950 1048 347006 1057
rect 346950 983 347006 992
rect 346964 480 346992 983
rect 348068 480 348096 2638
rect 348344 1193 348372 2774
rect 349402 2802 349430 3060
rect 350506 2825 350534 3060
rect 351610 2854 351638 3060
rect 351598 2848 351650 2854
rect 350492 2816 350548 2825
rect 349402 2774 349476 2802
rect 349250 2751 349306 2760
rect 348330 1184 348386 1193
rect 348330 1119 348386 1128
rect 349264 480 349292 2751
rect 349448 1057 349476 2774
rect 352714 2825 352742 3060
rect 353818 2961 353846 3060
rect 353804 2952 353860 2961
rect 353804 2887 353860 2896
rect 351598 2790 351650 2796
rect 352700 2816 352756 2825
rect 350492 2751 350548 2760
rect 354922 2802 354950 3060
rect 355048 2848 355100 2854
rect 354922 2774 354996 2802
rect 355048 2790 355100 2796
rect 356026 2802 356054 3060
rect 357130 2825 357158 3060
rect 358234 2854 358262 3060
rect 359338 2922 359366 3060
rect 360442 2961 360470 3060
rect 360428 2952 360484 2961
rect 359326 2916 359378 2922
rect 360428 2887 360484 2896
rect 359326 2858 359378 2864
rect 358222 2848 358274 2854
rect 356334 2816 356390 2825
rect 352700 2751 352756 2760
rect 353298 2680 353354 2689
rect 353354 2638 353616 2666
rect 353298 2615 353354 2624
rect 350446 1320 350502 1329
rect 350446 1255 350502 1264
rect 349434 1048 349490 1057
rect 349434 983 349490 992
rect 350460 480 350488 1255
rect 351642 1184 351698 1193
rect 351642 1119 351698 1128
rect 351656 480 351684 1119
rect 352838 1048 352894 1057
rect 352838 983 352894 992
rect 352852 480 352880 983
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 354 353616 2638
rect 354968 1329 354996 2774
rect 355060 1442 355088 2790
rect 356026 2774 356100 2802
rect 356072 2689 356100 2774
rect 356334 2751 356390 2760
rect 356886 2816 356942 2825
rect 357116 2816 357172 2825
rect 356942 2774 357020 2802
rect 356886 2751 356942 2760
rect 356058 2680 356114 2689
rect 356058 2615 356114 2624
rect 355060 1414 355272 1442
rect 354954 1320 355010 1329
rect 354954 1255 355010 1264
rect 355244 480 355272 1414
rect 356348 480 356376 2751
rect 356992 2666 357020 2774
rect 361546 2825 361574 3060
rect 361672 2848 361724 2854
rect 358222 2790 358274 2796
rect 359922 2816 359978 2825
rect 357116 2751 357172 2760
rect 359922 2751 359978 2760
rect 361118 2816 361174 2825
rect 361118 2751 361174 2760
rect 361532 2816 361588 2825
rect 362650 2802 362678 3060
rect 363754 2961 363782 3060
rect 363740 2952 363796 2961
rect 363328 2916 363380 2922
rect 363740 2887 363796 2896
rect 364064 2916 364116 2922
rect 363328 2858 363380 2864
rect 364064 2858 364116 2864
rect 361724 2796 361896 2802
rect 361672 2790 361896 2796
rect 361684 2774 361896 2790
rect 362650 2774 362724 2802
rect 361532 2751 361588 2760
rect 356992 2638 357572 2666
rect 357544 480 357572 2638
rect 358726 1320 358782 1329
rect 358726 1255 358782 1264
rect 358740 480 358768 1255
rect 359936 480 359964 2751
rect 361132 480 361160 2751
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 361868 354 361896 2774
rect 362696 1562 362724 2774
rect 363340 1578 363368 2858
rect 364076 2825 364104 2858
rect 364858 2825 364886 3060
rect 365962 2922 365990 3060
rect 365720 2916 365772 2922
rect 365720 2858 365772 2864
rect 365950 2916 366002 2922
rect 365950 2858 366002 2864
rect 364062 2816 364118 2825
rect 364062 2751 364118 2760
rect 364614 2816 364670 2825
rect 364614 2751 364670 2760
rect 364844 2816 364900 2825
rect 364844 2751 364900 2760
rect 362684 1556 362736 1562
rect 363340 1550 363552 1578
rect 362684 1498 362736 1504
rect 363524 480 363552 1550
rect 364628 480 364656 2751
rect 365732 1442 365760 2858
rect 367066 2854 367094 3060
rect 368170 2938 368198 3060
rect 368170 2910 368336 2938
rect 367054 2848 367106 2854
rect 367054 2790 367106 2796
rect 368202 2816 368258 2825
rect 368202 2751 368258 2760
rect 366824 1556 366876 1562
rect 366824 1498 366876 1504
rect 365732 1414 365852 1442
rect 365824 480 365852 1414
rect 366836 762 366864 1498
rect 366836 734 367048 762
rect 367020 480 367048 734
rect 368216 480 368244 2751
rect 368308 1562 368336 2910
rect 369274 2825 369302 3060
rect 370056 2922 370176 2938
rect 370378 2922 370406 3060
rect 370044 2916 370176 2922
rect 370096 2910 370176 2916
rect 370044 2858 370096 2864
rect 369260 2816 369316 2825
rect 369260 2751 369316 2760
rect 369030 2680 369086 2689
rect 369086 2638 369440 2666
rect 369030 2615 369086 2624
rect 368296 1556 368348 1562
rect 368296 1498 368348 1504
rect 369412 480 369440 2638
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370148 354 370176 2910
rect 370366 2916 370418 2922
rect 370366 2858 370418 2864
rect 371240 2848 371292 2854
rect 371332 2848 371384 2854
rect 371240 2790 371292 2796
rect 371330 2816 371332 2825
rect 371482 2825 371510 3060
rect 372586 2938 372614 3060
rect 373690 2961 373718 3060
rect 372540 2910 372614 2938
rect 373676 2952 373732 2961
rect 372540 2825 372568 2910
rect 373676 2887 373732 2896
rect 374000 2848 374052 2854
rect 371384 2816 371386 2825
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 2790
rect 371330 2751 371386 2760
rect 371468 2816 371524 2825
rect 371468 2751 371524 2760
rect 372526 2816 372582 2825
rect 374000 2790 374052 2796
rect 374794 2802 374822 3060
rect 375196 2916 375248 2922
rect 375196 2858 375248 2864
rect 372526 2751 372582 2760
rect 372620 1556 372672 1562
rect 372620 1498 372672 1504
rect 372632 1442 372660 1498
rect 374012 1442 374040 2790
rect 374794 2774 374868 2802
rect 374840 2689 374868 2774
rect 374826 2680 374882 2689
rect 374826 2615 374882 2624
rect 375208 1442 375236 2858
rect 375898 2854 375926 3060
rect 377002 2922 377030 3060
rect 376990 2916 377042 2922
rect 376990 2858 377042 2864
rect 375886 2848 375938 2854
rect 375886 2790 375938 2796
rect 376482 2816 376538 2825
rect 378106 2802 378134 3060
rect 379210 2825 379238 3060
rect 378874 2816 378930 2825
rect 378106 2786 378180 2802
rect 378106 2780 378192 2786
rect 378106 2774 378140 2780
rect 376482 2751 376538 2760
rect 372632 1414 372936 1442
rect 374012 1414 374132 1442
rect 375208 1414 375328 1442
rect 372908 480 372936 1414
rect 374104 480 374132 1414
rect 375300 480 375328 1414
rect 376496 480 376524 2751
rect 378874 2751 378930 2760
rect 379196 2816 379252 2825
rect 380314 2802 380342 3060
rect 380900 2848 380952 2854
rect 380314 2774 380388 2802
rect 381418 2825 381446 3060
rect 382522 2961 382550 3060
rect 382508 2952 382564 2961
rect 382280 2916 382332 2922
rect 382508 2887 382564 2896
rect 382280 2858 382332 2864
rect 380900 2790 380952 2796
rect 381404 2816 381460 2825
rect 379196 2751 379252 2760
rect 378140 2722 378192 2728
rect 377494 2544 377550 2553
rect 377550 2502 377720 2530
rect 377494 2479 377550 2488
rect 377692 480 377720 2502
rect 378888 480 378916 2751
rect 379518 2680 379574 2689
rect 379518 2615 379574 2624
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379532 354 379560 2615
rect 380360 1562 380388 2774
rect 380912 1578 380940 2790
rect 381404 2751 381460 2760
rect 382292 1578 382320 2858
rect 383626 2802 383654 3060
rect 384730 2904 384758 3060
rect 385834 2922 385862 3060
rect 385822 2916 385874 2922
rect 384730 2876 384988 2904
rect 384960 2825 384988 2876
rect 385822 2858 385874 2864
rect 383476 2780 383528 2786
rect 383476 2722 383528 2728
rect 383580 2774 383654 2802
rect 384762 2816 384818 2825
rect 383488 1578 383516 2722
rect 383580 2553 383608 2774
rect 384762 2751 384818 2760
rect 384946 2816 385002 2825
rect 386938 2802 386966 3060
rect 388042 2825 388070 3060
rect 389146 2854 389174 3060
rect 389134 2848 389186 2854
rect 387154 2816 387210 2825
rect 386938 2774 387012 2802
rect 384946 2751 385002 2760
rect 383566 2544 383622 2553
rect 383566 2479 383622 2488
rect 380348 1556 380400 1562
rect 380912 1550 381216 1578
rect 382292 1550 382412 1578
rect 383488 1550 383608 1578
rect 380348 1498 380400 1504
rect 381188 480 381216 1550
rect 382384 480 382412 1550
rect 383580 480 383608 1550
rect 384776 480 384804 2751
rect 386984 1562 387012 2774
rect 387154 2751 387210 2760
rect 387798 2816 387854 2825
rect 387798 2751 387854 2760
rect 388028 2816 388084 2825
rect 389134 2790 389186 2796
rect 390250 2802 390278 3060
rect 391354 2961 391382 3060
rect 392458 2961 392486 3060
rect 391340 2952 391396 2961
rect 392444 2952 392500 2961
rect 391340 2887 391396 2896
rect 391848 2916 391900 2922
rect 393562 2938 393590 3060
rect 392444 2887 392500 2896
rect 393228 2916 393280 2922
rect 391848 2858 391900 2864
rect 393562 2910 393636 2938
rect 394666 2922 394694 3060
rect 393228 2858 393280 2864
rect 390250 2774 390324 2802
rect 388028 2751 388084 2760
rect 385776 1556 385828 1562
rect 385776 1498 385828 1504
rect 386972 1556 387024 1562
rect 386972 1498 387024 1504
rect 385788 762 385816 1498
rect 385788 734 386000 762
rect 385972 480 386000 734
rect 387168 480 387196 2751
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 387812 354 387840 2751
rect 389454 2544 389510 2553
rect 389454 2479 389510 2488
rect 389468 480 389496 2479
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390296 105 390324 2774
rect 390558 2680 390614 2689
rect 390614 2638 390692 2666
rect 390558 2615 390614 2624
rect 390664 480 390692 2638
rect 391860 480 391888 2858
rect 393240 2825 393268 2858
rect 393504 2848 393556 2854
rect 393226 2816 393282 2825
rect 393226 2751 393282 2760
rect 393502 2816 393504 2825
rect 393556 2816 393558 2825
rect 393502 2751 393558 2760
rect 393608 1562 393636 2910
rect 394056 2916 394108 2922
rect 394654 2916 394706 2922
rect 394108 2876 394280 2904
rect 394056 2858 394108 2864
rect 392676 1556 392728 1562
rect 392676 1498 392728 1504
rect 393596 1556 393648 1562
rect 393596 1498 393648 1504
rect 390282 96 390338 105
rect 390282 31 390338 40
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392688 354 392716 1498
rect 394252 480 394280 2876
rect 394654 2858 394706 2864
rect 395770 2854 395798 3060
rect 395758 2848 395810 2854
rect 395342 2816 395398 2825
rect 396874 2825 396902 3060
rect 395758 2790 395810 2796
rect 396860 2816 396916 2825
rect 395342 2751 395398 2760
rect 397978 2802 398006 3060
rect 399082 2961 399110 3060
rect 399068 2952 399124 2961
rect 399068 2887 399124 2896
rect 400186 2802 400214 3060
rect 400864 2916 400916 2922
rect 400916 2876 401180 2904
rect 400864 2858 400916 2864
rect 397978 2774 398052 2802
rect 396860 2751 396916 2760
rect 395356 480 395384 2751
rect 397550 2680 397606 2689
rect 397606 2638 397776 2666
rect 397550 2615 397606 2624
rect 397748 480 397776 2638
rect 398024 1329 398052 2774
rect 400140 2774 400214 2802
rect 398838 2680 398894 2689
rect 398894 2638 398972 2666
rect 398838 2615 398894 2624
rect 398010 1320 398066 1329
rect 398010 1255 398066 1264
rect 398944 480 398972 2638
rect 399944 1556 399996 1562
rect 399944 1498 399996 1504
rect 399956 626 399984 1498
rect 400140 921 400168 2774
rect 401152 1578 401180 2876
rect 401290 2802 401318 3060
rect 402394 2961 402422 3060
rect 403498 2961 403526 3060
rect 402380 2952 402436 2961
rect 402380 2887 402436 2896
rect 403484 2952 403540 2961
rect 403484 2887 403540 2896
rect 404602 2854 404630 3060
rect 402336 2848 402388 2854
rect 401290 2774 401364 2802
rect 404590 2848 404642 2854
rect 402336 2790 402388 2796
rect 403622 2816 403678 2825
rect 401336 2009 401364 2774
rect 401322 2000 401378 2009
rect 401322 1935 401378 1944
rect 402348 1578 402376 2790
rect 405706 2802 405734 3060
rect 404590 2790 404642 2796
rect 403622 2751 403678 2760
rect 405660 2774 405734 2802
rect 406014 2816 406070 2825
rect 401152 1550 401364 1578
rect 402348 1550 402560 1578
rect 400126 912 400182 921
rect 400126 847 400182 856
rect 399956 598 400168 626
rect 400140 480 400168 598
rect 401336 480 401364 1550
rect 402532 480 402560 1550
rect 403636 480 403664 2751
rect 404818 1320 404874 1329
rect 404818 1255 404874 1264
rect 404832 480 404860 1255
rect 393014 354 393126 480
rect 392688 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396170 96 396226 105
rect 396510 82 396622 480
rect 396226 54 396622 82
rect 396170 31 396226 40
rect 396510 -960 396622 54
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405660 377 405688 2774
rect 406810 2802 406838 3060
rect 407914 2802 407942 3060
rect 409018 2961 409046 3060
rect 409004 2952 409060 2961
rect 409004 2887 409060 2896
rect 410122 2825 410150 3060
rect 409602 2816 409658 2825
rect 406810 2774 406884 2802
rect 407914 2774 407988 2802
rect 406014 2751 406070 2760
rect 406028 480 406056 2751
rect 406856 1329 406884 2774
rect 406842 1320 406898 1329
rect 406842 1255 406898 1264
rect 407210 640 407266 649
rect 407210 575 407266 584
rect 407224 480 407252 575
rect 405646 368 405702 377
rect 405646 303 405702 312
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 407960 105 407988 2774
rect 409602 2751 409658 2760
rect 410108 2816 410164 2825
rect 411226 2802 411254 3060
rect 410108 2751 410164 2760
rect 411180 2774 411254 2802
rect 411720 2848 411772 2854
rect 411720 2790 411772 2796
rect 412330 2802 412358 3060
rect 413434 2802 413462 3060
rect 414538 2802 414566 3060
rect 415642 2802 415670 3060
rect 416594 2816 416650 2825
rect 408406 2000 408462 2009
rect 408406 1935 408462 1944
rect 408420 480 408448 1935
rect 409616 480 409644 2751
rect 410430 2680 410486 2689
rect 410486 2638 410840 2666
rect 410430 2615 410486 2624
rect 410812 480 410840 2638
rect 411180 649 411208 2774
rect 411732 1578 411760 2790
rect 412330 2774 412404 2802
rect 413434 2774 413508 2802
rect 414538 2774 414612 2802
rect 415642 2774 415716 2802
rect 411732 1550 411944 1578
rect 411166 640 411222 649
rect 411166 575 411222 584
rect 411916 480 411944 1550
rect 412376 921 412404 2774
rect 413480 1057 413508 2774
rect 414294 1320 414350 1329
rect 414294 1255 414350 1264
rect 413466 1048 413522 1057
rect 413466 983 413522 992
rect 412362 912 412418 921
rect 412362 847 412418 856
rect 414308 480 414336 1255
rect 414584 513 414612 2774
rect 415688 1329 415716 2774
rect 416746 2802 416774 3060
rect 416594 2751 416650 2760
rect 416700 2774 416774 2802
rect 417850 2802 417878 3060
rect 417974 2816 418030 2825
rect 417850 2774 417924 2802
rect 415674 1320 415730 1329
rect 415674 1255 415730 1264
rect 416608 1034 416636 2751
rect 416700 1193 416728 2774
rect 416686 1184 416742 1193
rect 416686 1119 416742 1128
rect 416608 1006 416728 1034
rect 414570 504 414626 513
rect 407946 96 408002 105
rect 407946 31 408002 40
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412822 368 412878 377
rect 413070 354 413182 480
rect 412878 326 413182 354
rect 412822 303 412878 312
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 416700 480 416728 1006
rect 417896 785 417924 2774
rect 418954 2802 418982 3060
rect 420058 2802 420086 3060
rect 421162 2961 421190 3060
rect 421148 2952 421204 2961
rect 421148 2887 421204 2896
rect 422266 2802 422294 3060
rect 423370 2825 423398 3060
rect 418954 2774 419028 2802
rect 420058 2774 420132 2802
rect 417974 2751 418030 2760
rect 417882 776 417938 785
rect 417882 711 417938 720
rect 417988 626 418016 2751
rect 419000 2009 419028 2774
rect 418986 2000 419042 2009
rect 418986 1935 419042 1944
rect 420104 649 420132 2774
rect 422220 2774 422294 2802
rect 423356 2816 423412 2825
rect 421378 1048 421434 1057
rect 421378 983 421434 992
rect 420182 912 420238 921
rect 420182 847 420238 856
rect 417896 598 418016 626
rect 418986 640 419042 649
rect 417896 480 417924 598
rect 418986 575 419042 584
rect 420090 640 420146 649
rect 420090 575 420146 584
rect 419000 480 419028 575
rect 420196 480 420224 847
rect 421392 480 421420 983
rect 414570 439 414626 448
rect 415306 96 415362 105
rect 415462 82 415574 480
rect 415362 54 415574 82
rect 415306 31 415362 40
rect 415462 -960 415574 54
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422220 134 422248 2774
rect 424474 2802 424502 3060
rect 425578 2802 425606 3060
rect 426682 2802 426710 3060
rect 427786 2802 427814 3060
rect 424474 2774 424548 2802
rect 425578 2774 425652 2802
rect 426682 2774 426756 2802
rect 423356 2751 423412 2760
rect 424520 2145 424548 2774
rect 424506 2136 424562 2145
rect 424506 2071 424562 2080
rect 425624 1329 425652 2774
rect 423770 1320 423826 1329
rect 423770 1255 423826 1264
rect 425610 1320 425666 1329
rect 425610 1255 425666 1264
rect 423784 480 423812 1255
rect 424966 1184 425022 1193
rect 424966 1119 425022 1128
rect 424980 480 425008 1119
rect 426162 776 426218 785
rect 426162 711 426218 720
rect 426176 480 426204 711
rect 422546 354 422658 480
rect 422758 368 422814 377
rect 422546 326 422758 354
rect 422208 128 422260 134
rect 422208 70 422260 76
rect 422546 -960 422658 326
rect 422758 303 422814 312
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426728 241 426756 2774
rect 427740 2774 427814 2802
rect 428890 2802 428918 3060
rect 429994 2802 430022 3060
rect 431098 2802 431126 3060
rect 432050 2816 432106 2825
rect 428890 2774 428964 2802
rect 429994 2774 430068 2802
rect 431098 2774 431172 2802
rect 427740 2009 427768 2774
rect 427266 2000 427322 2009
rect 427266 1935 427322 1944
rect 427726 2000 427782 2009
rect 427726 1935 427782 1944
rect 427280 480 427308 1935
rect 428462 640 428518 649
rect 428462 575 428518 584
rect 428476 480 428504 575
rect 426714 232 426770 241
rect 426714 167 426770 176
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 428936 377 428964 2774
rect 429198 2680 429254 2689
rect 429198 2615 429254 2624
rect 428922 368 428978 377
rect 429212 354 429240 2615
rect 430040 2553 430068 2774
rect 430026 2544 430082 2553
rect 430026 2479 430082 2488
rect 431144 1358 431172 2774
rect 432202 2802 432230 3060
rect 433306 2802 433334 3060
rect 432202 2774 432276 2802
rect 432050 2751 432106 2760
rect 431132 1352 431184 1358
rect 431132 1294 431184 1300
rect 432064 480 432092 2751
rect 432248 1193 432276 2774
rect 433260 2774 433334 2802
rect 434410 2802 434438 3060
rect 435514 2802 435542 3060
rect 436618 2802 436646 3060
rect 437722 2802 437750 3060
rect 438826 2802 438854 3060
rect 434410 2774 434484 2802
rect 435514 2774 435588 2802
rect 436618 2774 436692 2802
rect 437722 2774 437796 2802
rect 433260 2417 433288 2774
rect 433246 2408 433302 2417
rect 433246 2343 433302 2352
rect 433246 2136 433302 2145
rect 433246 2071 433302 2080
rect 432234 1184 432290 1193
rect 432234 1119 432290 1128
rect 433260 480 433288 2071
rect 434456 1737 434484 2774
rect 435560 2281 435588 2774
rect 435546 2272 435602 2281
rect 435546 2207 435602 2216
rect 436664 2145 436692 2774
rect 436650 2136 436706 2145
rect 436650 2071 436706 2080
rect 437768 2009 437796 2774
rect 438780 2774 438854 2802
rect 439930 2802 439958 3060
rect 441034 2802 441062 3060
rect 442138 2802 442166 3060
rect 443242 2802 443270 3060
rect 444346 2802 444374 3060
rect 439930 2774 440004 2802
rect 441034 2774 441108 2802
rect 442138 2774 442212 2802
rect 443242 2774 443316 2802
rect 436742 2000 436798 2009
rect 436742 1935 436798 1944
rect 437754 2000 437810 2009
rect 437754 1935 437810 1944
rect 434442 1728 434498 1737
rect 434442 1663 434498 1672
rect 434442 1320 434498 1329
rect 434442 1255 434498 1264
rect 434456 480 434484 1255
rect 435376 598 435588 626
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 428922 303 428978 312
rect 429630 -960 429742 326
rect 430826 82 430938 480
rect 431040 128 431092 134
rect 430826 76 431040 82
rect 430826 70 431092 76
rect 430826 54 431080 70
rect 430826 -960 430938 54
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435376 241 435404 598
rect 435560 480 435588 598
rect 436756 480 436784 1935
rect 435362 232 435418 241
rect 435362 167 435418 176
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437478 368 437534 377
rect 437910 354 438022 480
rect 437534 326 438022 354
rect 437478 303 437534 312
rect 437910 -960 438022 326
rect 438780 202 438808 2774
rect 439134 2544 439190 2553
rect 439134 2479 439190 2488
rect 439148 480 439176 2479
rect 439976 1873 440004 2774
rect 441080 2689 441108 2774
rect 441066 2680 441122 2689
rect 441066 2615 441122 2624
rect 442184 2553 442212 2774
rect 442170 2544 442226 2553
rect 442170 2479 442226 2488
rect 443288 2417 443316 2774
rect 444300 2774 444374 2802
rect 445450 2802 445478 3060
rect 446554 2802 446582 3060
rect 447658 2802 447686 3060
rect 448762 2802 448790 3060
rect 449866 2854 449894 3060
rect 449854 2848 449906 2854
rect 445450 2774 445524 2802
rect 446554 2774 446628 2802
rect 447658 2774 447732 2802
rect 448762 2774 448836 2802
rect 449854 2790 449906 2796
rect 450970 2802 450998 3060
rect 452074 2961 452102 3060
rect 453178 2961 453206 3060
rect 452060 2952 452116 2961
rect 452060 2887 452116 2896
rect 453164 2952 453220 2961
rect 453164 2887 453220 2896
rect 454282 2802 454310 3060
rect 455386 2961 455414 3060
rect 456490 2961 456518 3060
rect 455372 2952 455428 2961
rect 455372 2887 455428 2896
rect 456476 2952 456532 2961
rect 456476 2887 456532 2896
rect 450970 2774 451044 2802
rect 454282 2774 454356 2802
rect 442630 2408 442686 2417
rect 442630 2343 442686 2352
rect 443274 2408 443330 2417
rect 443274 2343 443330 2352
rect 439962 1864 440018 1873
rect 439962 1799 440018 1808
rect 439964 1352 440016 1358
rect 439964 1294 440016 1300
rect 438768 196 438820 202
rect 438768 138 438820 144
rect 439106 -960 439218 480
rect 439976 218 440004 1294
rect 441526 1184 441582 1193
rect 441526 1119 441582 1128
rect 441540 480 441568 1119
rect 442644 480 442672 2343
rect 443826 1728 443882 1737
rect 443826 1663 443882 1672
rect 443840 480 443868 1663
rect 440302 218 440414 480
rect 439976 190 440414 218
rect 440302 -960 440414 190
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444300 134 444328 2774
rect 445496 2281 445524 2774
rect 445022 2272 445078 2281
rect 445022 2207 445078 2216
rect 445482 2272 445538 2281
rect 445482 2207 445538 2216
rect 445036 480 445064 2207
rect 446600 2145 446628 2774
rect 446218 2136 446274 2145
rect 446218 2071 446274 2080
rect 446586 2136 446642 2145
rect 446586 2071 446642 2080
rect 446232 480 446260 2071
rect 447414 2000 447470 2009
rect 447414 1935 447470 1944
rect 447428 480 447456 1935
rect 447704 513 447732 2774
rect 448808 2009 448836 2774
rect 450910 2680 450966 2689
rect 450910 2615 450966 2624
rect 448794 2000 448850 2009
rect 448794 1935 448850 1944
rect 449806 1864 449862 1873
rect 449806 1799 449862 1808
rect 447690 504 447746 513
rect 444288 128 444340 134
rect 444288 70 444340 76
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 449820 480 449848 1799
rect 450924 480 450952 2615
rect 451016 1358 451044 2774
rect 452106 2544 452162 2553
rect 452106 2479 452162 2488
rect 451004 1352 451056 1358
rect 451004 1294 451056 1300
rect 452120 480 452148 2479
rect 453302 2408 453358 2417
rect 453302 2343 453358 2352
rect 453316 480 453344 2343
rect 454328 1290 454356 2774
rect 457594 2774 457622 3060
rect 458698 2961 458726 3060
rect 459802 2961 459830 3060
rect 458684 2952 458740 2961
rect 458684 2887 458740 2896
rect 459788 2952 459844 2961
rect 459788 2887 459844 2896
rect 460388 2848 460440 2854
rect 460388 2790 460440 2796
rect 457594 2746 457668 2774
rect 455694 2272 455750 2281
rect 455694 2207 455750 2216
rect 454316 1284 454368 1290
rect 454316 1226 454368 1232
rect 455708 480 455736 2207
rect 456890 2136 456946 2145
rect 456890 2071 456946 2080
rect 456904 480 456932 2071
rect 447690 439 447746 448
rect 448582 218 448694 480
rect 448440 202 448694 218
rect 448428 196 448694 202
rect 448480 190 448694 196
rect 448428 138 448480 144
rect 448582 -960 448694 190
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454132 128 454184 134
rect 454470 82 454582 480
rect 454184 76 454582 82
rect 454132 70 454582 76
rect 454144 54 454582 70
rect 454470 -960 454582 54
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 457640 105 457668 2746
rect 459190 2000 459246 2009
rect 459190 1935 459246 1944
rect 457916 598 458128 626
rect 457718 504 457774 513
rect 457916 490 457944 598
rect 457774 462 457944 490
rect 458100 480 458128 598
rect 459204 480 459232 1935
rect 460400 480 460428 2790
rect 460906 2774 460934 3060
rect 460860 2746 460934 2774
rect 462010 2774 462038 3060
rect 463114 2774 463142 3060
rect 464218 2961 464246 3060
rect 464204 2952 464260 2961
rect 464204 2887 464260 2896
rect 463974 2816 464030 2825
rect 462010 2746 462084 2774
rect 463114 2746 463188 2774
rect 463974 2751 464030 2760
rect 465322 2774 465350 3060
rect 466426 2774 466454 3060
rect 467530 2802 467558 3060
rect 468634 2802 468662 3060
rect 469738 2802 469766 3060
rect 470842 2938 470870 3060
rect 471946 2961 471974 3060
rect 471932 2952 471988 2961
rect 470842 2910 471284 2938
rect 471256 2825 471284 2910
rect 471932 2887 471988 2896
rect 469862 2816 469918 2825
rect 467530 2774 467604 2802
rect 468634 2774 468708 2802
rect 469738 2774 469812 2802
rect 457718 439 457774 448
rect 457626 96 457682 105
rect 457626 31 457682 40
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 460860 134 460888 2746
rect 462056 1358 462084 2746
rect 462686 2680 462742 2689
rect 462742 2638 462820 2666
rect 462686 2615 462742 2624
rect 461308 1352 461360 1358
rect 461308 1294 461360 1300
rect 462044 1352 462096 1358
rect 462044 1294 462096 1300
rect 461320 762 461348 1294
rect 461320 734 461624 762
rect 461596 480 461624 734
rect 462792 480 462820 2638
rect 463160 2281 463188 2746
rect 463146 2272 463202 2281
rect 463146 2207 463202 2216
rect 463988 480 464016 2751
rect 465322 2746 465396 2774
rect 465080 1284 465132 1290
rect 465132 1244 465212 1272
rect 465080 1226 465132 1232
rect 465184 480 465212 1244
rect 465368 513 465396 2746
rect 466380 2746 466454 2774
rect 466274 2544 466330 2553
rect 466274 2479 466330 2488
rect 465354 504 465410 513
rect 460848 128 460900 134
rect 460848 70 460900 76
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466288 480 466316 2479
rect 466380 1222 466408 2746
rect 467286 2544 467342 2553
rect 467342 2502 467512 2530
rect 467286 2479 467342 2488
rect 466368 1216 466420 1222
rect 466368 1158 466420 1164
rect 467484 480 467512 2502
rect 467576 1358 467604 2774
rect 468680 2145 468708 2774
rect 468666 2136 468722 2145
rect 468666 2071 468722 2080
rect 469784 2009 469812 2774
rect 469862 2751 469918 2760
rect 471058 2816 471114 2825
rect 471058 2751 471114 2760
rect 471242 2816 471298 2825
rect 473050 2802 473078 3060
rect 474154 2802 474182 3060
rect 475258 2802 475286 3060
rect 476362 2802 476390 3060
rect 477466 2802 477494 3060
rect 473050 2774 473124 2802
rect 474154 2774 474228 2802
rect 475258 2774 475332 2802
rect 471242 2751 471298 2760
rect 469770 2000 469826 2009
rect 469770 1935 469826 1944
rect 467564 1352 467616 1358
rect 467564 1294 467616 1300
rect 468496 598 468708 626
rect 465354 439 465410 448
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468496 105 468524 598
rect 468680 480 468708 598
rect 469876 480 469904 2751
rect 471072 480 471100 2751
rect 473096 1358 473124 2774
rect 472992 1352 473044 1358
rect 472992 1294 473044 1300
rect 473084 1352 473136 1358
rect 473084 1294 473136 1300
rect 473004 1154 473032 1294
rect 473360 1284 473412 1290
rect 473360 1226 473412 1232
rect 472992 1148 473044 1154
rect 472992 1090 473044 1096
rect 473372 626 473400 1226
rect 473372 598 473492 626
rect 473464 480 473492 598
rect 468482 96 468538 105
rect 468482 31 468538 40
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 82 472338 480
rect 472440 128 472492 134
rect 472226 76 472440 82
rect 472226 70 472492 76
rect 472226 54 472480 70
rect 472226 -960 472338 54
rect 473422 -960 473534 480
rect 474200 202 474228 2774
rect 474554 2272 474610 2281
rect 474554 2207 474610 2216
rect 474568 480 474596 2207
rect 475304 785 475332 2774
rect 476316 2774 476390 2802
rect 477420 2774 477494 2802
rect 478570 2802 478598 3060
rect 478880 2848 478932 2854
rect 478570 2774 478644 2802
rect 478880 2790 478932 2796
rect 479674 2802 479702 3060
rect 480778 2802 480806 3060
rect 481882 2802 481910 3060
rect 482834 2816 482890 2825
rect 475382 2680 475438 2689
rect 475438 2638 475792 2666
rect 475382 2615 475438 2624
rect 475290 776 475346 785
rect 475290 711 475346 720
rect 475764 480 475792 2638
rect 474188 196 474240 202
rect 474188 138 474240 144
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476316 105 476344 2774
rect 476394 504 476450 513
rect 476450 462 476528 490
rect 476394 439 476450 448
rect 476500 354 476528 462
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476302 96 476358 105
rect 476302 31 476358 40
rect 476918 -960 477030 326
rect 477420 134 477448 2774
rect 477868 1216 477920 1222
rect 477868 1158 477920 1164
rect 477880 626 477908 1158
rect 477880 598 478184 626
rect 478156 480 478184 598
rect 478616 513 478644 2774
rect 478892 1358 478920 2790
rect 479674 2774 479748 2802
rect 480778 2774 480852 2802
rect 481882 2774 481956 2802
rect 479720 1358 479748 2774
rect 480534 2136 480590 2145
rect 480534 2071 480590 2080
rect 478880 1352 478932 1358
rect 478880 1294 478932 1300
rect 479708 1352 479760 1358
rect 479708 1294 479760 1300
rect 478892 1154 479012 1170
rect 478880 1148 479012 1154
rect 478932 1142 479012 1148
rect 478880 1090 478932 1096
rect 478602 504 478658 513
rect 477408 128 477460 134
rect 477408 70 477460 76
rect 478114 -960 478226 480
rect 478602 439 478658 448
rect 478984 354 479012 1142
rect 480548 480 480576 2071
rect 480824 649 480852 2774
rect 481730 2000 481786 2009
rect 481730 1935 481786 1944
rect 480810 640 480866 649
rect 480810 575 480866 584
rect 481744 480 481772 1935
rect 481928 921 481956 2774
rect 482986 2802 483014 3060
rect 482834 2751 482890 2760
rect 482940 2774 483014 2802
rect 483938 2816 483994 2825
rect 481914 912 481970 921
rect 481914 847 481970 856
rect 482848 480 482876 2751
rect 482940 678 482968 2774
rect 484090 2802 484118 3060
rect 485194 2961 485222 3060
rect 485180 2952 485236 2961
rect 485180 2887 485236 2896
rect 485228 2848 485280 2854
rect 484090 2774 484256 2802
rect 486298 2802 486326 3060
rect 487402 2802 487430 3060
rect 488506 2802 488534 3060
rect 485228 2790 485280 2796
rect 483938 2751 483994 2760
rect 483952 1986 483980 2751
rect 483952 1958 484072 1986
rect 482928 672 482980 678
rect 482928 614 482980 620
rect 484044 480 484072 1958
rect 479310 354 479422 480
rect 478984 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484228 270 484256 2774
rect 485240 480 485268 2790
rect 486160 2774 486326 2802
rect 487264 2774 487430 2802
rect 488460 2774 488534 2802
rect 489610 2802 489638 3060
rect 490714 2802 490742 3060
rect 491818 2825 491846 3060
rect 489610 2774 489684 2802
rect 484216 264 484268 270
rect 484216 206 484268 212
rect 485198 -960 485310 480
rect 486160 377 486188 2774
rect 486146 368 486202 377
rect 486146 303 486202 312
rect 486394 218 486506 480
rect 487264 241 487292 2774
rect 488460 1290 488488 2774
rect 488448 1284 488500 1290
rect 488448 1226 488500 1232
rect 487618 776 487674 785
rect 487618 711 487674 720
rect 487632 480 487660 711
rect 487250 232 487306 241
rect 486394 202 486648 218
rect 486394 196 486660 202
rect 486394 190 486608 196
rect 486394 -960 486506 190
rect 487250 167 487306 176
rect 486608 138 486660 144
rect 487590 -960 487702 480
rect 488786 82 488898 480
rect 489656 105 489684 2774
rect 490668 2774 490742 2802
rect 491804 2816 491860 2825
rect 488998 96 489054 105
rect 488786 54 488998 82
rect 488786 -960 488898 54
rect 488998 31 489054 40
rect 489642 96 489698 105
rect 489642 31 489698 40
rect 489890 82 490002 480
rect 490668 202 490696 2774
rect 492922 2802 492950 3060
rect 494026 2802 494054 3060
rect 495130 2961 495158 3060
rect 495116 2952 495172 2961
rect 495116 2887 495172 2896
rect 492922 2774 492996 2802
rect 491804 2751 491860 2760
rect 492036 1352 492088 1358
rect 492036 1294 492088 1300
rect 492048 762 492076 1294
rect 492048 734 492352 762
rect 490746 504 490802 513
rect 492324 480 492352 734
rect 492968 513 492996 2774
rect 493980 2774 494054 2802
rect 496234 2802 496262 3060
rect 497338 2802 497366 3060
rect 498442 2802 498470 3060
rect 499546 2802 499574 3060
rect 496234 2774 496308 2802
rect 497338 2774 497412 2802
rect 498442 2774 498516 2802
rect 493506 640 493562 649
rect 493506 575 493562 584
rect 492954 504 493010 513
rect 490746 439 490802 448
rect 490760 354 490788 439
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 490656 196 490708 202
rect 490656 138 490708 144
rect 490104 128 490156 134
rect 489890 76 490104 82
rect 489890 70 490156 76
rect 489890 54 490144 70
rect 489890 -960 490002 54
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493520 480 493548 575
rect 492954 439 493010 448
rect 493478 -960 493590 480
rect 493980 134 494008 2774
rect 496280 1358 496308 2774
rect 496268 1352 496320 1358
rect 496268 1294 496320 1300
rect 494702 912 494758 921
rect 494702 847 494758 856
rect 494716 480 494744 847
rect 497384 746 497412 2774
rect 498198 2544 498254 2553
rect 498198 2479 498254 2488
rect 497372 740 497424 746
rect 497372 682 497424 688
rect 495900 672 495952 678
rect 495900 614 495952 620
rect 495912 480 495940 614
rect 498212 480 498240 2479
rect 498488 649 498516 2774
rect 499500 2774 499574 2802
rect 500650 2802 500678 3060
rect 501754 2802 501782 3060
rect 502858 2802 502886 3060
rect 503962 2802 503990 3060
rect 505066 2802 505094 3060
rect 500650 2774 500724 2802
rect 501754 2774 502104 2802
rect 499500 678 499528 2774
rect 500696 814 500724 2774
rect 501696 1284 501748 1290
rect 501696 1226 501748 1232
rect 500684 808 500736 814
rect 500684 750 500736 756
rect 499488 672 499540 678
rect 498474 640 498530 649
rect 501708 660 501736 1226
rect 501708 632 501828 660
rect 499488 614 499540 620
rect 498474 575 498530 584
rect 500328 598 500632 626
rect 493968 128 494020 134
rect 493968 70 494020 76
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 218 497178 480
rect 497280 264 497332 270
rect 497066 212 497280 218
rect 497066 206 497332 212
rect 497066 190 497320 206
rect 497066 -960 497178 190
rect 498170 -960 498282 480
rect 498934 368 498990 377
rect 499366 354 499478 480
rect 498990 326 499478 354
rect 498934 303 498990 312
rect 499366 -960 499478 326
rect 500328 241 500356 598
rect 500604 480 500632 598
rect 501800 480 501828 632
rect 500314 232 500370 241
rect 500314 167 500370 176
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502076 377 502104 2774
rect 502720 2774 502886 2802
rect 503732 2774 503990 2802
rect 505020 2774 505094 2802
rect 505374 2816 505430 2825
rect 502062 368 502118 377
rect 502062 303 502118 312
rect 502720 241 502748 2774
rect 502706 232 502762 241
rect 502706 167 502762 176
rect 502954 82 503066 480
rect 503732 105 503760 2774
rect 504150 218 504262 480
rect 505020 270 505048 2774
rect 506170 2802 506198 3060
rect 507274 2802 507302 3060
rect 508378 2961 508406 3060
rect 508364 2952 508420 2961
rect 508364 2887 508420 2896
rect 509482 2825 509510 3060
rect 506170 2774 506244 2802
rect 505374 2751 505430 2760
rect 505388 480 505416 2751
rect 503824 202 504262 218
rect 505008 264 505060 270
rect 505008 206 505060 212
rect 503812 196 504262 202
rect 503864 190 504262 196
rect 503812 138 503864 144
rect 503166 96 503222 105
rect 502954 54 503166 82
rect 502954 -960 503066 54
rect 503166 31 503222 40
rect 503718 96 503774 105
rect 503718 31 503774 40
rect 504150 -960 504262 190
rect 505346 -960 505458 480
rect 506216 406 506244 2774
rect 507228 2774 507302 2802
rect 508870 2816 508926 2825
rect 506662 504 506718 513
rect 506204 400 506256 406
rect 506204 342 506256 348
rect 506450 354 506562 480
rect 506662 439 506718 448
rect 506676 354 506704 439
rect 506450 326 506704 354
rect 506450 -960 506562 326
rect 507228 202 507256 2774
rect 508870 2751 508926 2760
rect 509468 2816 509524 2825
rect 510586 2802 510614 3060
rect 511690 2961 511718 3060
rect 511676 2952 511732 2961
rect 511676 2887 511732 2896
rect 512794 2825 512822 3060
rect 509468 2751 509524 2760
rect 510540 2774 510614 2802
rect 512780 2816 512836 2825
rect 508884 480 508912 2751
rect 509608 1352 509660 1358
rect 509608 1294 509660 1300
rect 507216 196 507268 202
rect 507216 138 507268 144
rect 507308 128 507360 134
rect 507646 82 507758 480
rect 507360 76 507758 82
rect 507308 70 507758 76
rect 507320 54 507758 70
rect 507646 -960 507758 54
rect 508842 -960 508954 480
rect 509620 354 509648 1294
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 510540 134 510568 2774
rect 513898 2802 513926 3060
rect 515002 2961 515030 3060
rect 514988 2952 515044 2961
rect 514988 2887 515044 2896
rect 516106 2802 516134 3060
rect 513898 2774 513972 2802
rect 512780 2751 512836 2760
rect 513944 746 513972 2774
rect 516060 2774 516134 2802
rect 517210 2802 517238 3060
rect 518314 2961 518342 3060
rect 518300 2952 518356 2961
rect 518300 2887 518356 2896
rect 519418 2802 519446 3060
rect 517210 2774 517376 2802
rect 516060 1290 516088 2774
rect 516048 1284 516100 1290
rect 516048 1226 516100 1232
rect 514760 808 514812 814
rect 514760 750 514812 756
rect 513932 740 513984 746
rect 513932 682 513984 688
rect 512458 640 512514 649
rect 512458 575 512514 584
rect 512472 480 512500 575
rect 514772 480 514800 750
rect 517150 640 517206 649
rect 517150 575 517206 584
rect 517164 480 517192 575
rect 511234 354 511346 480
rect 511448 468 511500 474
rect 511448 410 511500 416
rect 511460 354 511488 410
rect 511234 326 511488 354
rect 510528 128 510580 134
rect 510528 70 510580 76
rect 511234 -960 511346 326
rect 512430 -960 512542 480
rect 513534 354 513646 480
rect 513392 338 513646 354
rect 513380 332 513646 338
rect 513432 326 513646 332
rect 513380 274 513432 280
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515494 368 515550 377
rect 515926 354 516038 480
rect 515550 326 516038 354
rect 515494 303 515550 312
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517348 338 517376 2774
rect 519372 2774 519446 2802
rect 520522 2802 520550 3060
rect 521626 2802 521654 3060
rect 520522 2774 520596 2802
rect 518176 598 518388 626
rect 517336 332 517388 338
rect 517336 274 517388 280
rect 518176 105 518204 598
rect 518360 480 518388 598
rect 519372 513 519400 2774
rect 519358 504 519414 513
rect 518162 96 518218 105
rect 518162 31 518218 40
rect 518318 -960 518430 480
rect 519358 439 519414 448
rect 519514 218 519626 480
rect 520568 270 520596 2774
rect 521580 2774 521654 2802
rect 522730 2802 522758 3060
rect 523834 2802 523862 3060
rect 524938 2961 524966 3060
rect 524924 2952 524980 2961
rect 524924 2887 524980 2896
rect 524234 2816 524290 2825
rect 522730 2774 522804 2802
rect 523834 2774 523908 2802
rect 521580 1154 521608 2774
rect 521568 1148 521620 1154
rect 521568 1090 521620 1096
rect 520740 672 520792 678
rect 520740 614 520792 620
rect 520752 480 520780 614
rect 519728 264 519780 270
rect 519514 212 519728 218
rect 519514 206 519780 212
rect 520556 264 520608 270
rect 520556 206 520608 212
rect 519514 190 519768 206
rect 519514 -960 519626 190
rect 520710 -960 520822 480
rect 521814 218 521926 480
rect 521672 202 521926 218
rect 522776 202 522804 2774
rect 523038 2544 523094 2553
rect 523038 2479 523094 2488
rect 523052 480 523080 2479
rect 521660 196 521926 202
rect 521712 190 521926 196
rect 521660 138 521712 144
rect 521814 -960 521926 190
rect 522764 196 522816 202
rect 522764 138 522816 144
rect 523010 -960 523122 480
rect 523880 406 523908 2774
rect 524234 2751 524290 2760
rect 526042 2774 526070 3060
rect 527146 2774 527174 3060
rect 524248 480 524276 2751
rect 526042 2746 526116 2774
rect 523868 400 523920 406
rect 523868 342 523920 348
rect 524206 -960 524318 480
rect 525402 82 525514 480
rect 526088 241 526116 2746
rect 527100 2746 527174 2774
rect 528250 2774 528278 3060
rect 529354 2961 529382 3060
rect 529340 2952 529396 2961
rect 529340 2887 529396 2896
rect 530458 2774 530486 3060
rect 531562 2961 531590 3060
rect 531548 2952 531604 2961
rect 531548 2887 531604 2896
rect 532666 2774 532694 3060
rect 528250 2746 528324 2774
rect 530458 2746 530532 2774
rect 526534 2680 526590 2689
rect 526590 2638 526668 2666
rect 526534 2615 526590 2624
rect 526640 480 526668 2638
rect 526074 232 526130 241
rect 526074 167 526130 176
rect 525616 128 525668 134
rect 525402 76 525616 82
rect 525402 70 525668 76
rect 525402 54 525656 70
rect 525402 -960 525514 54
rect 526598 -960 526710 480
rect 527100 134 527128 2746
rect 527638 2680 527694 2689
rect 527694 2638 527864 2666
rect 527638 2615 527694 2624
rect 527836 480 527864 2638
rect 528296 2009 528324 2746
rect 530030 2680 530086 2689
rect 530086 2638 530164 2666
rect 530030 2615 530086 2624
rect 528282 2000 528338 2009
rect 528282 1935 528338 1944
rect 529020 740 529072 746
rect 529020 682 529072 688
rect 529032 480 529060 682
rect 530136 480 530164 2638
rect 530504 1222 530532 2746
rect 532620 2746 532694 2774
rect 533770 2774 533798 3060
rect 534874 2802 534902 3060
rect 535978 2961 536006 3060
rect 535964 2952 536020 2961
rect 535964 2887 536020 2896
rect 537082 2802 537110 3060
rect 538186 2802 538214 3060
rect 534874 2774 534948 2802
rect 537082 2774 537156 2802
rect 533770 2746 533844 2774
rect 531320 1284 531372 1290
rect 531320 1226 531372 1232
rect 530492 1216 530544 1222
rect 530492 1158 530544 1164
rect 531332 480 531360 1226
rect 532620 626 532648 2746
rect 533342 2680 533398 2689
rect 533398 2638 533752 2666
rect 533342 2615 533398 2624
rect 532620 598 532740 626
rect 527088 128 527140 134
rect 527088 70 527140 76
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 354 532598 480
rect 532160 338 532598 354
rect 532712 338 532740 598
rect 533724 480 533752 2638
rect 533816 1358 533844 2746
rect 533804 1352 533856 1358
rect 533804 1294 533856 1300
rect 534920 785 534948 2774
rect 537128 1290 537156 2774
rect 538140 2774 538214 2802
rect 539290 2802 539318 3060
rect 540394 2802 540422 3060
rect 541498 2961 541526 3060
rect 541484 2952 541540 2961
rect 541484 2887 541540 2896
rect 542602 2825 542630 3060
rect 540794 2816 540850 2825
rect 539290 2774 539364 2802
rect 540394 2774 540468 2802
rect 537116 1284 537168 1290
rect 537116 1226 537168 1232
rect 537036 1154 537248 1170
rect 537024 1148 537248 1154
rect 537076 1142 537248 1148
rect 537024 1090 537076 1096
rect 534906 776 534962 785
rect 534906 711 534962 720
rect 534736 598 534948 626
rect 532148 332 532598 338
rect 532200 326 532598 332
rect 532148 274 532200 280
rect 532486 -960 532598 326
rect 532700 332 532752 338
rect 532700 274 532752 280
rect 533682 -960 533794 480
rect 534736 105 534764 598
rect 534920 480 534948 598
rect 537220 480 537248 1142
rect 534722 96 534778 105
rect 534722 31 534778 40
rect 534878 -960 534990 480
rect 536074 218 536186 480
rect 536288 264 536340 270
rect 536074 212 536288 218
rect 536074 206 536340 212
rect 536074 190 536328 206
rect 536074 -960 536186 190
rect 537178 -960 537290 480
rect 538140 270 538168 2774
rect 538128 264 538180 270
rect 538374 218 538486 480
rect 539336 474 539364 2774
rect 539324 468 539376 474
rect 539324 410 539376 416
rect 538128 206 538180 212
rect 538232 202 538486 218
rect 538220 196 538486 202
rect 538272 190 538486 196
rect 538220 138 538272 144
rect 538374 -960 538486 190
rect 539570 354 539682 480
rect 539784 400 539836 406
rect 539570 348 539784 354
rect 539570 342 539836 348
rect 539570 326 539824 342
rect 539570 -960 539682 326
rect 540440 202 540468 2774
rect 540794 2751 540850 2760
rect 542588 2816 542644 2825
rect 543706 2802 543734 3060
rect 542588 2751 542644 2760
rect 543660 2774 543734 2802
rect 544810 2774 544838 3060
rect 545914 2774 545942 3060
rect 547018 2774 547046 3060
rect 548122 2961 548150 3060
rect 548108 2952 548164 2961
rect 548108 2887 548164 2896
rect 549226 2774 549254 3060
rect 540808 480 540836 2751
rect 540428 196 540480 202
rect 540428 138 540480 144
rect 540766 -960 540878 480
rect 541962 218 542074 480
rect 542174 232 542230 241
rect 541962 190 542174 218
rect 541962 -960 542074 190
rect 542174 167 542230 176
rect 542820 128 542872 134
rect 543158 82 543270 480
rect 543660 134 543688 2774
rect 544810 2746 544884 2774
rect 545914 2746 545988 2774
rect 547018 2746 547092 2774
rect 544382 2000 544438 2009
rect 544382 1935 544438 1944
rect 544396 480 544424 1935
rect 542872 76 543270 82
rect 542820 70 543270 76
rect 543648 128 543700 134
rect 543648 70 543700 76
rect 542832 54 543270 70
rect 543158 -960 543270 54
rect 544354 -960 544466 480
rect 544856 105 544884 2746
rect 545302 2544 545358 2553
rect 545358 2502 545528 2530
rect 545302 2479 545358 2488
rect 545500 480 545528 2502
rect 545960 785 545988 2746
rect 546500 1216 546552 1222
rect 546500 1158 546552 1164
rect 545946 776 546002 785
rect 545946 711 546002 720
rect 544842 96 544898 105
rect 544842 31 544898 40
rect 545458 -960 545570 480
rect 546512 354 546540 1158
rect 546654 354 546766 480
rect 547064 406 547092 2746
rect 549180 2746 549254 2774
rect 550330 2774 550358 3060
rect 551434 2774 551462 3060
rect 550330 2746 550404 2774
rect 547878 2544 547934 2553
rect 547878 2479 547934 2488
rect 547892 480 547920 2479
rect 549180 1154 549208 2746
rect 550088 1352 550140 1358
rect 550088 1294 550140 1300
rect 549168 1148 549220 1154
rect 549168 1090 549220 1096
rect 550100 762 550128 1294
rect 550376 1290 550404 2746
rect 551388 2746 551462 2774
rect 552538 2774 552566 3060
rect 553642 2802 553670 3060
rect 554746 2802 554774 3060
rect 553642 2774 553716 2802
rect 552538 2746 552612 2774
rect 550364 1284 550416 1290
rect 550364 1226 550416 1232
rect 550100 734 550312 762
rect 550284 480 550312 734
rect 551388 649 551416 2746
rect 552478 2680 552534 2689
rect 552478 2615 552534 2624
rect 552492 762 552520 2615
rect 552584 921 552612 2746
rect 553688 1358 553716 2774
rect 554700 2774 554774 2802
rect 555850 2802 555878 3060
rect 556954 2802 556982 3060
rect 555850 2774 555924 2802
rect 553676 1352 553728 1358
rect 553676 1294 553728 1300
rect 553768 1216 553820 1222
rect 553768 1158 553820 1164
rect 552570 912 552626 921
rect 552570 847 552626 856
rect 552492 734 552704 762
rect 551374 640 551430 649
rect 551374 575 551430 584
rect 551480 598 551692 626
rect 551480 480 551508 598
rect 546512 326 546766 354
rect 547052 400 547104 406
rect 547052 342 547104 348
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 549046 354 549158 480
rect 548720 338 549158 354
rect 548708 332 549158 338
rect 548760 326 549158 332
rect 548708 274 548760 280
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 551664 377 551692 598
rect 552676 480 552704 734
rect 553780 480 553808 1158
rect 551650 368 551706 377
rect 551650 303 551706 312
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554700 338 554728 2774
rect 555896 1222 555924 2774
rect 556908 2774 556982 2802
rect 558058 2802 558086 3060
rect 558550 2816 558606 2825
rect 558058 2774 558132 2802
rect 555884 1216 555936 1222
rect 555884 1158 555936 1164
rect 554688 332 554740 338
rect 554688 274 554740 280
rect 554780 264 554832 270
rect 554934 218 555046 480
rect 554832 212 555046 218
rect 554780 206 555046 212
rect 554792 190 555046 206
rect 554934 -960 555046 190
rect 556130 354 556242 480
rect 556344 468 556396 474
rect 556344 410 556396 416
rect 556356 354 556384 410
rect 556130 326 556384 354
rect 556130 -960 556242 326
rect 556908 270 556936 2774
rect 556896 264 556948 270
rect 557326 218 557438 480
rect 558104 377 558132 2774
rect 559162 2802 559190 3060
rect 560266 2802 560294 3060
rect 559162 2774 559236 2802
rect 558550 2751 558606 2760
rect 558564 480 558592 2751
rect 559208 513 559236 2774
rect 560220 2774 560294 2802
rect 561370 2802 561398 3060
rect 562474 2802 562502 3060
rect 563578 2802 563606 3060
rect 565634 2816 565690 2825
rect 561370 2774 561444 2802
rect 562474 2774 562548 2802
rect 563578 2774 563652 2802
rect 559286 2544 559342 2553
rect 559342 2502 559420 2530
rect 559286 2479 559342 2488
rect 559194 504 559250 513
rect 558090 368 558146 377
rect 558090 303 558146 312
rect 556896 206 556948 212
rect 557000 202 557438 218
rect 556988 196 557438 202
rect 557040 190 557438 196
rect 556988 138 557040 144
rect 557326 -960 557438 190
rect 558522 -960 558634 480
rect 559194 439 559250 448
rect 559392 354 559420 2502
rect 559718 354 559830 480
rect 559392 326 559830 354
rect 559718 -960 559830 326
rect 560220 202 560248 2774
rect 560208 196 560260 202
rect 560208 138 560260 144
rect 560484 128 560536 134
rect 560822 82 560934 480
rect 561416 134 561444 2774
rect 560536 76 560934 82
rect 560484 70 560934 76
rect 561404 128 561456 134
rect 561404 70 561456 76
rect 562018 82 562130 480
rect 562520 241 562548 2774
rect 563242 776 563298 785
rect 563242 711 563298 720
rect 563256 480 563284 711
rect 562506 232 562562 241
rect 562506 167 562562 176
rect 562230 96 562286 105
rect 560496 54 560934 70
rect 560822 -960 560934 54
rect 562018 54 562230 82
rect 562018 -960 562130 54
rect 562230 31 562286 40
rect 563214 -960 563326 480
rect 563624 105 563652 2774
rect 565634 2751 565690 2760
rect 565648 480 565676 2751
rect 571064 1352 571116 1358
rect 571064 1294 571116 1300
rect 567568 1284 567620 1290
rect 567568 1226 567620 1232
rect 566832 1148 566884 1154
rect 566832 1090 566884 1096
rect 566844 480 566872 1090
rect 564410 354 564522 480
rect 564624 400 564676 406
rect 564410 348 564624 354
rect 564410 342 564676 348
rect 564410 326 564664 342
rect 563610 96 563666 105
rect 563610 31 563666 40
rect 564410 -960 564522 326
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567580 354 567608 1226
rect 570326 912 570382 921
rect 570326 847 570382 856
rect 569130 640 569186 649
rect 569130 575 569186 584
rect 569144 480 569172 575
rect 570340 480 570368 847
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571076 354 571104 1294
rect 573364 1216 573416 1222
rect 573364 1158 573416 1164
rect 571494 354 571606 480
rect 571076 326 571606 354
rect 571494 -960 571606 326
rect 572690 354 572802 480
rect 573376 354 573404 1158
rect 577134 504 577190 513
rect 573886 354 573998 480
rect 572690 338 572944 354
rect 572690 332 572956 338
rect 572690 326 572904 332
rect 572690 -960 572802 326
rect 573376 326 573998 354
rect 572904 274 572956 280
rect 573886 -960 573998 326
rect 575082 218 575194 480
rect 575754 368 575810 377
rect 576278 354 576390 480
rect 577134 439 577190 448
rect 575810 326 576390 354
rect 577148 354 577176 439
rect 577382 354 577494 480
rect 577148 326 577494 354
rect 575754 303 575810 312
rect 575296 264 575348 270
rect 575082 212 575296 218
rect 575082 206 575348 212
rect 575082 190 575336 206
rect 575082 -960 575194 190
rect 576278 -960 576390 326
rect 577382 -960 577494 326
rect 578578 218 578690 480
rect 578578 202 578832 218
rect 578578 196 578844 202
rect 578578 190 578792 196
rect 578578 -960 578690 190
rect 578792 138 578844 144
rect 579774 -960 579886 480
rect 580970 82 581082 480
rect 581826 232 581882 241
rect 582166 218 582278 480
rect 581882 190 582278 218
rect 581826 167 581882 176
rect 581184 128 581236 134
rect 580970 76 581184 82
rect 580970 70 581236 76
rect 580970 54 581224 70
rect 580970 -960 581082 54
rect 582166 -960 582278 190
rect 583362 82 583474 480
rect 583574 96 583630 105
rect 583362 54 583574 82
rect 583362 -960 583474 54
rect 583574 31 583630 40
<< via2 >>
rect 17038 2760 17094 2816
rect 6458 992 6514 1048
rect 5262 856 5318 912
rect 4066 584 4122 640
rect 8758 720 8814 776
rect 386 40 442 96
rect 1490 176 1546 232
rect 3330 312 3386 368
rect 8206 448 8262 504
rect 10966 992 11022 1048
rect 12346 992 12402 1048
rect 11702 856 11758 912
rect 9586 584 9642 640
rect 11150 584 11206 640
rect 19246 1028 19248 1048
rect 19248 1028 19300 1048
rect 19300 1028 19302 1048
rect 19246 992 19302 1028
rect 19430 856 19486 912
rect 17866 720 17922 776
rect 18234 720 18290 776
rect 20350 40 20406 96
rect 21822 992 21878 1048
rect 21454 176 21510 232
rect 23018 2760 23074 2816
rect 23846 992 23902 1048
rect 22558 312 22614 368
rect 24766 312 24822 368
rect 28262 584 28318 640
rect 26330 176 26386 232
rect 26974 448 27030 504
rect 28170 448 28226 504
rect 35852 2896 35908 2952
rect 31022 856 31078 912
rect 31298 584 31354 640
rect 30286 312 30342 368
rect 33230 584 33286 640
rect 34794 2488 34850 2544
rect 36910 720 36966 776
rect 37002 448 37058 504
rect 41372 2760 41428 2816
rect 40774 2624 40830 2680
rect 44638 176 44694 232
rect 44638 40 44694 96
rect 47858 2624 47914 2680
rect 52412 2896 52468 2952
rect 53010 2624 53066 2680
rect 57932 2760 57988 2816
rect 58438 2760 58494 2816
rect 59634 1944 59690 2000
rect 64326 2760 64382 2816
rect 68972 2896 69028 2952
rect 65522 2080 65578 2136
rect 61198 40 61254 96
rect 66994 2216 67050 2272
rect 74492 2896 74548 2952
rect 69110 2352 69166 2408
rect 72606 2488 72662 2544
rect 76194 2760 76250 2816
rect 75550 1944 75606 2000
rect 77390 584 77446 640
rect 81070 2080 81126 2136
rect 82174 2216 82230 2272
rect 84382 2352 84438 2408
rect 83462 448 83518 504
rect 84658 312 84714 368
rect 87694 2488 87750 2544
rect 87786 312 87842 368
rect 91052 2760 91108 2816
rect 91558 2760 91614 2816
rect 92110 584 92166 640
rect 90178 40 90234 96
rect 93950 1944 94006 2000
rect 97630 448 97686 504
rect 99746 2216 99802 2272
rect 98826 448 98882 504
rect 101034 2080 101090 2136
rect 102230 2352 102286 2408
rect 102046 720 102102 776
rect 105404 2760 105460 2816
rect 105726 2488 105782 2544
rect 104162 40 104218 96
rect 107566 1944 107622 2000
rect 108118 1944 108174 2000
rect 109314 2624 109370 2680
rect 111614 1808 111670 1864
rect 113086 2216 113142 2272
rect 115294 2352 115350 2408
rect 114190 2080 114246 2136
rect 115202 2080 115258 2136
rect 112810 1672 112866 1728
rect 117686 2760 117742 2816
rect 118606 2488 118662 2544
rect 121918 2624 121974 2680
rect 120814 1944 120870 2000
rect 124126 1808 124182 1864
rect 125230 1672 125286 1728
rect 123482 720 123538 776
rect 119158 40 119214 96
rect 125690 176 125746 232
rect 127438 2080 127494 2136
rect 129692 2760 129748 2816
rect 129370 856 129426 912
rect 130566 584 130622 640
rect 132774 992 132830 1048
rect 127162 312 127218 368
rect 130750 448 130806 504
rect 132774 584 132830 640
rect 132958 584 133014 640
rect 135258 1944 135314 2000
rect 135166 720 135222 776
rect 136454 720 136510 776
rect 137282 176 137338 232
rect 137466 176 137522 232
rect 138478 312 138534 368
rect 141238 2216 141294 2272
rect 140686 856 140742 912
rect 142434 2080 142490 2136
rect 141790 992 141846 1048
rect 143538 2352 143594 2408
rect 147126 2760 147182 2816
rect 146206 1944 146262 2000
rect 143998 584 144054 640
rect 148322 1944 148378 2000
rect 147310 720 147366 776
rect 139858 40 139914 96
rect 148506 448 148562 504
rect 149518 2488 149574 2544
rect 150346 40 150402 96
rect 150622 2624 150678 2680
rect 151726 2216 151782 2272
rect 152830 2080 152886 2136
rect 151818 1808 151874 1864
rect 153934 2352 153990 2408
rect 154210 2080 154266 2136
rect 155406 2216 155462 2272
rect 157292 2760 157348 2816
rect 156602 2352 156658 2408
rect 160558 2624 160614 2680
rect 159454 2488 159510 2544
rect 158350 1944 158406 2000
rect 161294 1944 161350 2000
rect 157798 1672 157854 1728
rect 159270 40 159326 96
rect 160282 448 160338 504
rect 162490 2488 162546 2544
rect 161662 1808 161718 1864
rect 166078 2352 166134 2408
rect 164974 2216 165030 2272
rect 163870 2080 163926 2136
rect 167182 1672 167238 1728
rect 164882 1264 164938 1320
rect 167182 720 167238 776
rect 165894 312 165950 368
rect 168378 992 168434 1048
rect 168010 40 168066 96
rect 169390 448 169446 504
rect 171598 2488 171654 2544
rect 170494 1944 170550 2000
rect 173806 1264 173862 1320
rect 174266 1264 174322 1320
rect 171966 1128 172022 1184
rect 170586 448 170642 504
rect 173162 584 173218 640
rect 177118 992 177174 1048
rect 177854 992 177910 1048
rect 176014 720 176070 776
rect 174910 312 174966 368
rect 175830 40 175886 96
rect 179050 720 179106 776
rect 180246 1944 180302 2000
rect 176842 312 176898 368
rect 179326 448 179382 504
rect 180430 1128 180486 1184
rect 181442 856 181498 912
rect 182638 1264 182694 1320
rect 181534 584 181590 640
rect 182362 176 182418 232
rect 183466 40 183522 96
rect 183742 1128 183798 1184
rect 184938 1264 184994 1320
rect 184846 584 184902 640
rect 186134 2760 186190 2816
rect 185950 992 186006 1048
rect 188158 1944 188214 2000
rect 189722 1944 189778 2000
rect 189262 856 189318 912
rect 187054 720 187110 776
rect 187146 40 187202 96
rect 188986 312 189042 368
rect 193724 2760 193780 2816
rect 192574 1264 192630 1320
rect 191470 1128 191526 1184
rect 194414 1128 194470 1184
rect 193218 992 193274 1048
rect 192022 856 192078 912
rect 190826 720 190882 776
rect 190366 176 190422 232
rect 195610 1264 195666 1320
rect 196990 1944 197046 2000
rect 200302 992 200358 1048
rect 199198 856 199254 912
rect 200486 1672 200542 1728
rect 201498 1400 201554 1456
rect 201406 1128 201462 1184
rect 198094 720 198150 776
rect 199106 720 199162 776
rect 195886 584 195942 640
rect 202510 1264 202566 1320
rect 202694 992 202750 1048
rect 194782 40 194838 96
rect 197174 40 197230 96
rect 198370 312 198426 368
rect 203890 1128 203946 1184
rect 203522 40 203578 96
rect 205086 1264 205142 1320
rect 207386 2080 207442 2136
rect 206926 1672 206982 1728
rect 206190 1536 206246 1592
rect 205822 720 205878 776
rect 208582 1944 208638 2000
rect 208030 1400 208086 1456
rect 209778 2216 209834 2272
rect 209134 992 209190 1048
rect 212170 1808 212226 1864
rect 211342 1264 211398 1320
rect 210238 1128 210294 1184
rect 210974 1128 211030 1184
rect 213550 2080 213606 2136
rect 216862 2352 216918 2408
rect 215758 2216 215814 2272
rect 214654 1944 214710 2000
rect 213366 1672 213422 1728
rect 212446 1536 212502 1592
rect 215666 1536 215722 1592
rect 214470 1400 214526 1456
rect 218058 2624 218114 2680
rect 217966 1808 218022 1864
rect 216954 1128 217010 1184
rect 219254 2216 219310 2272
rect 219070 1672 219126 1728
rect 220450 1944 220506 2000
rect 220174 1400 220230 1456
rect 223486 2624 223542 2680
rect 222382 2352 222438 2408
rect 224590 2216 224646 2272
rect 223946 2080 224002 2136
rect 221554 1808 221610 1864
rect 221278 1536 221334 1592
rect 222750 1672 222806 1728
rect 225694 1944 225750 2000
rect 227534 1944 227590 2000
rect 226798 1808 226854 1864
rect 226338 1536 226394 1592
rect 225142 1400 225198 1456
rect 228730 2352 228786 2408
rect 227902 1672 227958 1728
rect 229006 2080 229062 2136
rect 229834 2080 229890 2136
rect 233422 2352 233478 2408
rect 234526 2080 234582 2136
rect 232318 1944 232374 2000
rect 233422 1808 233478 1864
rect 231214 1536 231270 1592
rect 232226 1536 232282 1592
rect 230110 1400 230166 1456
rect 231030 1400 231086 1456
rect 234618 1672 234674 1728
rect 238114 1944 238170 2000
rect 237838 1808 237894 1864
rect 236734 1536 236790 1592
rect 237010 1536 237066 1592
rect 235630 1400 235686 1456
rect 235814 1400 235870 1456
rect 239310 2080 239366 2136
rect 238942 1672 238998 1728
rect 243358 2080 243414 2136
rect 242254 1944 242310 2000
rect 241702 1808 241758 1864
rect 241150 1536 241206 1592
rect 240046 1400 240102 1456
rect 240506 1400 240562 1456
rect 242898 1672 242954 1728
rect 244094 1536 244150 1592
rect 246394 2352 246450 2408
rect 245566 1808 245622 1864
rect 244462 1400 244518 1456
rect 245198 1400 245254 1456
rect 247590 1808 247646 1864
rect 246670 1672 246726 1728
rect 248786 1944 248842 2000
rect 247774 1536 247830 1592
rect 249982 2352 250038 2408
rect 252190 1944 252246 2000
rect 251086 1808 251142 1864
rect 251178 1672 251234 1728
rect 249982 1536 250038 1592
rect 248878 1400 248934 1456
rect 254398 1672 254454 1728
rect 254674 1672 254730 1728
rect 253294 1536 253350 1592
rect 253478 1536 253534 1592
rect 252374 1400 252430 1456
rect 257710 1672 257766 1728
rect 258262 1672 258318 1728
rect 256606 1536 256662 1592
rect 257066 1536 257122 1592
rect 255502 1400 255558 1456
rect 255870 1400 255926 1456
rect 261022 1672 261078 1728
rect 261758 1672 261814 1728
rect 259918 1536 259974 1592
rect 260654 1536 260710 1592
rect 258814 1400 258870 1456
rect 259458 1264 259514 1320
rect 264334 1672 264390 1728
rect 263230 1536 263286 1592
rect 264150 1536 264206 1592
rect 262954 1400 263010 1456
rect 262126 1264 262182 1320
rect 266542 1536 266598 1592
rect 265438 1400 265494 1456
rect 266542 1128 266598 1184
rect 265346 992 265402 1048
rect 267738 1264 267794 1320
rect 267646 992 267702 1048
rect 268842 1400 268898 1456
rect 268750 1128 268806 1184
rect 270038 1536 270094 1592
rect 269854 1264 269910 1320
rect 272062 1536 272118 1592
rect 270958 1400 271014 1456
rect 271234 1264 271290 1320
rect 273166 1264 273222 1320
rect 273626 1264 273682 1320
rect 272430 1128 272486 1184
rect 275374 1264 275430 1320
rect 276018 1264 276074 1320
rect 274270 1128 274326 1184
rect 274822 1128 274878 1184
rect 277582 1264 277638 1320
rect 279514 1264 279570 1320
rect 276478 1128 276534 1184
rect 277122 1128 277178 1184
rect 278686 1128 278742 1184
rect 278318 992 278374 1048
rect 280894 1264 280950 1320
rect 281906 1264 281962 1320
rect 280710 1128 280766 1184
rect 279790 992 279846 1048
rect 283194 1264 283250 1320
rect 281998 1128 282054 1184
rect 285402 1264 285458 1320
rect 286414 1264 286470 1320
rect 286598 1264 286654 1320
rect 287518 1264 287574 1320
rect 287794 1264 287850 1320
rect 288622 1264 288678 1320
rect 204718 312 204774 368
rect 313002 1264 313058 1320
rect 313830 1264 313886 1320
rect 314106 1264 314162 1320
rect 315026 1264 315082 1320
rect 315210 1264 315266 1320
rect 316222 1264 316278 1320
rect 317418 1264 317474 1320
rect 318522 1264 318578 1320
rect 319626 1264 319682 1320
rect 318430 1128 318486 1184
rect 320914 1264 320970 1320
rect 319718 1128 319774 1184
rect 320730 1128 320786 1184
rect 322846 1264 322902 1320
rect 324410 1264 324466 1320
rect 325146 1264 325202 1320
rect 322110 1128 322166 1184
rect 324042 1128 324098 1184
rect 321834 992 321890 1048
rect 323306 992 323362 1048
rect 326802 1264 326858 1320
rect 327354 1264 327410 1320
rect 325606 1128 325662 1184
rect 326250 1128 326306 1184
rect 329194 1264 329250 1320
rect 329562 1264 329618 1320
rect 327998 1128 328054 1184
rect 328366 1128 328422 1184
rect 331586 1264 331642 1320
rect 330390 1128 330446 1184
rect 330666 1128 330722 1184
rect 332690 1128 332746 1184
rect 332874 1128 332930 1184
rect 331770 856 331826 912
rect 335082 1264 335138 1320
rect 335082 1128 335138 1184
rect 336186 1128 336242 1184
rect 333886 992 333942 1048
rect 333886 856 333942 912
rect 337474 1264 337530 1320
rect 338394 1264 338450 1320
rect 336278 992 336334 1048
rect 337290 992 337346 1048
rect 338670 1128 338726 1184
rect 339406 1128 339462 1184
rect 340970 1264 341026 1320
rect 341706 1264 341762 1320
rect 339866 992 339922 1048
rect 340602 992 340658 1048
rect 342166 1128 342222 1184
rect 342810 1128 342866 1184
rect 344972 2760 345028 2816
rect 346076 2760 346132 2816
rect 347778 2624 347834 2680
rect 344558 1264 344614 1320
rect 347226 1264 347282 1320
rect 343362 992 343418 1048
rect 343914 992 343970 1048
rect 345754 1128 345810 1184
rect 346950 992 347006 1048
rect 349250 2760 349306 2816
rect 348330 1128 348386 1184
rect 350492 2760 350548 2816
rect 353804 2896 353860 2952
rect 352700 2760 352756 2816
rect 360428 2896 360484 2952
rect 353298 2624 353354 2680
rect 350446 1264 350502 1320
rect 349434 992 349490 1048
rect 351642 1128 351698 1184
rect 352838 992 352894 1048
rect 356334 2760 356390 2816
rect 356886 2760 356942 2816
rect 356058 2624 356114 2680
rect 354954 1264 355010 1320
rect 357116 2760 357172 2816
rect 359922 2760 359978 2816
rect 361118 2760 361174 2816
rect 361532 2760 361588 2816
rect 363740 2896 363796 2952
rect 358726 1264 358782 1320
rect 364062 2760 364118 2816
rect 364614 2760 364670 2816
rect 364844 2760 364900 2816
rect 368202 2760 368258 2816
rect 369260 2760 369316 2816
rect 369030 2624 369086 2680
rect 373676 2896 373732 2952
rect 371330 2796 371332 2816
rect 371332 2796 371384 2816
rect 371384 2796 371386 2816
rect 371330 2760 371386 2796
rect 371468 2760 371524 2816
rect 372526 2760 372582 2816
rect 374826 2624 374882 2680
rect 376482 2760 376538 2816
rect 378874 2760 378930 2816
rect 379196 2760 379252 2816
rect 382508 2896 382564 2952
rect 377494 2488 377550 2544
rect 379518 2624 379574 2680
rect 381404 2760 381460 2816
rect 384762 2760 384818 2816
rect 384946 2760 385002 2816
rect 383566 2488 383622 2544
rect 387154 2760 387210 2816
rect 387798 2760 387854 2816
rect 388028 2760 388084 2816
rect 391340 2896 391396 2952
rect 392444 2896 392500 2952
rect 389454 2488 389510 2544
rect 390558 2624 390614 2680
rect 393226 2760 393282 2816
rect 393502 2796 393504 2816
rect 393504 2796 393556 2816
rect 393556 2796 393558 2816
rect 393502 2760 393558 2796
rect 390282 40 390338 96
rect 395342 2760 395398 2816
rect 396860 2760 396916 2816
rect 399068 2896 399124 2952
rect 397550 2624 397606 2680
rect 398838 2624 398894 2680
rect 398010 1264 398066 1320
rect 402380 2896 402436 2952
rect 403484 2896 403540 2952
rect 401322 1944 401378 2000
rect 403622 2760 403678 2816
rect 400126 856 400182 912
rect 404818 1264 404874 1320
rect 396170 40 396226 96
rect 406014 2760 406070 2816
rect 409004 2896 409060 2952
rect 406842 1264 406898 1320
rect 407210 584 407266 640
rect 405646 312 405702 368
rect 409602 2760 409658 2816
rect 410108 2760 410164 2816
rect 408406 1944 408462 2000
rect 410430 2624 410486 2680
rect 411166 584 411222 640
rect 414294 1264 414350 1320
rect 413466 992 413522 1048
rect 412362 856 412418 912
rect 416594 2760 416650 2816
rect 415674 1264 415730 1320
rect 416686 1128 416742 1184
rect 407946 40 408002 96
rect 412822 312 412878 368
rect 414570 448 414626 504
rect 417974 2760 418030 2816
rect 421148 2896 421204 2952
rect 417882 720 417938 776
rect 418986 1944 419042 2000
rect 421378 992 421434 1048
rect 420182 856 420238 912
rect 418986 584 419042 640
rect 420090 584 420146 640
rect 415306 40 415362 96
rect 423356 2760 423412 2816
rect 424506 2080 424562 2136
rect 423770 1264 423826 1320
rect 425610 1264 425666 1320
rect 424966 1128 425022 1184
rect 426162 720 426218 776
rect 422758 312 422814 368
rect 427266 1944 427322 2000
rect 427726 1944 427782 2000
rect 428462 584 428518 640
rect 426714 176 426770 232
rect 429198 2624 429254 2680
rect 428922 312 428978 368
rect 430026 2488 430082 2544
rect 432050 2760 432106 2816
rect 433246 2352 433302 2408
rect 433246 2080 433302 2136
rect 432234 1128 432290 1184
rect 435546 2216 435602 2272
rect 436650 2080 436706 2136
rect 436742 1944 436798 2000
rect 437754 1944 437810 2000
rect 434442 1672 434498 1728
rect 434442 1264 434498 1320
rect 435362 176 435418 232
rect 437478 312 437534 368
rect 439134 2488 439190 2544
rect 441066 2624 441122 2680
rect 442170 2488 442226 2544
rect 452060 2896 452116 2952
rect 453164 2896 453220 2952
rect 455372 2896 455428 2952
rect 456476 2896 456532 2952
rect 442630 2352 442686 2408
rect 443274 2352 443330 2408
rect 439962 1808 440018 1864
rect 441526 1128 441582 1184
rect 443826 1672 443882 1728
rect 445022 2216 445078 2272
rect 445482 2216 445538 2272
rect 446218 2080 446274 2136
rect 446586 2080 446642 2136
rect 447414 1944 447470 2000
rect 450910 2624 450966 2680
rect 448794 1944 448850 2000
rect 449806 1808 449862 1864
rect 447690 448 447746 504
rect 452106 2488 452162 2544
rect 453302 2352 453358 2408
rect 458684 2896 458740 2952
rect 459788 2896 459844 2952
rect 455694 2216 455750 2272
rect 456890 2080 456946 2136
rect 459190 1944 459246 2000
rect 457718 448 457774 504
rect 464204 2896 464260 2952
rect 463974 2760 464030 2816
rect 471932 2896 471988 2952
rect 457626 40 457682 96
rect 462686 2624 462742 2680
rect 463146 2216 463202 2272
rect 466274 2488 466330 2544
rect 465354 448 465410 504
rect 467286 2488 467342 2544
rect 468666 2080 468722 2136
rect 469862 2760 469918 2816
rect 471058 2760 471114 2816
rect 471242 2760 471298 2816
rect 469770 1944 469826 2000
rect 468482 40 468538 96
rect 474554 2216 474610 2272
rect 475382 2624 475438 2680
rect 475290 720 475346 776
rect 476394 448 476450 504
rect 476302 40 476358 96
rect 480534 2080 480590 2136
rect 478602 448 478658 504
rect 481730 1944 481786 2000
rect 480810 584 480866 640
rect 482834 2760 482890 2816
rect 481914 856 481970 912
rect 483938 2760 483994 2816
rect 485180 2896 485236 2952
rect 486146 312 486202 368
rect 487618 720 487674 776
rect 487250 176 487306 232
rect 488998 40 489054 96
rect 489642 40 489698 96
rect 491804 2760 491860 2816
rect 495116 2896 495172 2952
rect 490746 448 490802 504
rect 493506 584 493562 640
rect 492954 448 493010 504
rect 494702 856 494758 912
rect 498198 2488 498254 2544
rect 498474 584 498530 640
rect 498934 312 498990 368
rect 500314 176 500370 232
rect 502062 312 502118 368
rect 502706 176 502762 232
rect 505374 2760 505430 2816
rect 508364 2896 508420 2952
rect 503166 40 503222 96
rect 503718 40 503774 96
rect 506662 448 506718 504
rect 508870 2760 508926 2816
rect 509468 2760 509524 2816
rect 511676 2896 511732 2952
rect 512780 2760 512836 2816
rect 514988 2896 515044 2952
rect 518300 2896 518356 2952
rect 512458 584 512514 640
rect 517150 584 517206 640
rect 515494 312 515550 368
rect 518162 40 518218 96
rect 519358 448 519414 504
rect 524924 2896 524980 2952
rect 523038 2488 523094 2544
rect 524234 2760 524290 2816
rect 529340 2896 529396 2952
rect 531548 2896 531604 2952
rect 526534 2624 526590 2680
rect 526074 176 526130 232
rect 527638 2624 527694 2680
rect 530030 2624 530086 2680
rect 528282 1944 528338 2000
rect 535964 2896 536020 2952
rect 533342 2624 533398 2680
rect 541484 2896 541540 2952
rect 534906 720 534962 776
rect 534722 40 534778 96
rect 540794 2760 540850 2816
rect 542588 2760 542644 2816
rect 548108 2896 548164 2952
rect 542174 176 542230 232
rect 544382 1944 544438 2000
rect 545302 2488 545358 2544
rect 545946 720 546002 776
rect 544842 40 544898 96
rect 547878 2488 547934 2544
rect 552478 2624 552534 2680
rect 552570 856 552626 912
rect 551374 584 551430 640
rect 551650 312 551706 368
rect 558550 2760 558606 2816
rect 559286 2488 559342 2544
rect 558090 312 558146 368
rect 559194 448 559250 504
rect 563242 720 563298 776
rect 562506 176 562562 232
rect 562230 40 562286 96
rect 565634 2760 565690 2816
rect 563610 40 563666 96
rect 570326 856 570382 912
rect 569130 584 569186 640
rect 575754 312 575810 368
rect 577134 448 577190 504
rect 581826 176 581882 232
rect 583574 40 583630 96
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371378 480 371468
rect 3734 371378 3740 371380
rect -960 371318 3740 371378
rect -960 371228 480 371318
rect 3734 371316 3740 371318
rect 3804 371316 3810 371380
rect 583520 364972 584960 365212
rect -960 358458 480 358548
rect 3550 358458 3556 358460
rect -960 358398 3556 358458
rect -960 358308 480 358398
rect 3550 358396 3556 358398
rect 3620 358396 3626 358460
rect 583520 351780 584960 352020
rect -960 345402 480 345492
rect 3366 345402 3372 345404
rect -960 345342 3372 345402
rect -960 345252 480 345342
rect 3366 345340 3372 345342
rect 3436 345340 3442 345404
rect 3734 344660 3740 344724
rect 3804 344722 3810 344724
rect 574686 344722 574692 344724
rect 3804 344662 12052 344722
rect 571964 344662 574692 344722
rect 3804 344660 3810 344662
rect 574686 344660 574692 344662
rect 574756 344660 574762 344724
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 3550 330244 3556 330308
rect 3620 330306 3626 330308
rect 574870 330306 574876 330308
rect 3620 330246 12052 330306
rect 571964 330246 574876 330306
rect 3620 330244 3626 330246
rect 574870 330244 574876 330246
rect 574940 330244 574946 330308
rect 574686 325212 574692 325276
rect 574756 325274 574762 325276
rect 583520 325274 584960 325364
rect 574756 325214 584960 325274
rect 574756 325212 574762 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3734 319290 3740 319292
rect -960 319230 3740 319290
rect -960 319140 480 319230
rect 3734 319228 3740 319230
rect 3804 319228 3810 319292
rect 3366 315828 3372 315892
rect 3436 315890 3442 315892
rect 575054 315890 575060 315892
rect 3436 315830 12052 315890
rect 571964 315830 575060 315890
rect 3436 315828 3442 315830
rect 575054 315828 575060 315830
rect 575124 315828 575130 315892
rect 574870 312020 574876 312084
rect 574940 312082 574946 312084
rect 583520 312082 584960 312172
rect 574940 312022 584960 312082
rect 574940 312020 574946 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3550 306234 3556 306236
rect -960 306174 3556 306234
rect -960 306084 480 306174
rect 3550 306172 3556 306174
rect 3620 306172 3626 306236
rect 3734 301412 3740 301476
rect 3804 301474 3810 301476
rect 574686 301474 574692 301476
rect 3804 301414 12052 301474
rect 571964 301414 574692 301474
rect 3804 301412 3810 301414
rect 574686 301412 574692 301414
rect 574756 301412 574762 301476
rect 575054 298692 575060 298756
rect 575124 298754 575130 298756
rect 583520 298754 584960 298844
rect 575124 298694 584960 298754
rect 575124 298692 575130 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3366 293178 3372 293180
rect -960 293118 3372 293178
rect -960 293028 480 293118
rect 3366 293116 3372 293118
rect 3436 293116 3442 293180
rect 3550 286996 3556 287060
rect 3620 287058 3626 287060
rect 575054 287058 575060 287060
rect 3620 286998 12052 287058
rect 571964 286998 575060 287058
rect 3620 286996 3626 286998
rect 575054 286996 575060 286998
rect 575124 286996 575130 287060
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 3366 272580 3372 272644
rect 3436 272642 3442 272644
rect 574870 272642 574876 272644
rect 3436 272582 12052 272642
rect 571964 272582 574876 272642
rect 3436 272580 3442 272582
rect 574870 272580 574876 272582
rect 574940 272580 574946 272644
rect 574686 272172 574692 272236
rect 574756 272234 574762 272236
rect 583520 272234 584960 272324
rect 574756 272174 584960 272234
rect 574756 272172 574762 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 8150 267202 8156 267204
rect -960 267142 8156 267202
rect -960 267052 480 267142
rect 8150 267140 8156 267142
rect 8220 267140 8226 267204
rect 575054 258844 575060 258908
rect 575124 258906 575130 258908
rect 583520 258906 584960 258996
rect 575124 258846 584960 258906
rect 575124 258844 575130 258846
rect 583520 258756 584960 258846
rect 8150 258164 8156 258228
rect 8220 258226 8226 258228
rect 574686 258226 574692 258228
rect 8220 258166 12052 258226
rect 571964 258166 574692 258226
rect 8220 258164 8226 258166
rect 574686 258164 574692 258166
rect 574756 258164 574762 258228
rect -960 254146 480 254236
rect 7414 254146 7420 254148
rect -960 254086 7420 254146
rect -960 253996 480 254086
rect 7414 254084 7420 254086
rect 7484 254084 7490 254148
rect 574870 245516 574876 245580
rect 574940 245578 574946 245580
rect 583520 245578 584960 245668
rect 574940 245518 584960 245578
rect 574940 245516 574946 245518
rect 583520 245428 584960 245518
rect 7414 243748 7420 243812
rect 7484 243810 7490 243812
rect 574870 243810 574876 243812
rect 7484 243750 12052 243810
rect 571964 243750 574876 243810
rect 7484 243748 7490 243750
rect 574870 243748 574876 243750
rect 574940 243748 574946 243812
rect -960 241090 480 241180
rect 7414 241090 7420 241092
rect -960 241030 7420 241090
rect -960 240940 480 241030
rect 7414 241028 7420 241030
rect 7484 241028 7490 241092
rect 574686 232324 574692 232388
rect 574756 232386 574762 232388
rect 583520 232386 584960 232476
rect 574756 232326 584960 232386
rect 574756 232324 574762 232326
rect 583520 232236 584960 232326
rect 7414 229332 7420 229396
rect 7484 229394 7490 229396
rect 574686 229394 574692 229396
rect 7484 229334 12052 229394
rect 571964 229334 574692 229394
rect 7484 229332 7490 229334
rect 574686 229332 574692 229334
rect 574756 229332 574762 229396
rect -960 227884 480 228124
rect 574870 218996 574876 219060
rect 574940 219058 574946 219060
rect 583520 219058 584960 219148
rect 574940 218998 584960 219058
rect 574940 218996 574946 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 574870 214978 574876 214980
rect -960 214918 12052 214978
rect 571964 214918 574876 214978
rect -960 214828 480 214918
rect 574870 214916 574876 214918
rect 574940 214916 574946 214980
rect 574686 205668 574692 205732
rect 574756 205730 574762 205732
rect 583520 205730 584960 205820
rect 574756 205670 584960 205730
rect 574756 205668 574762 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect -960 201862 6930 201922
rect -960 201772 480 201862
rect 6870 201242 6930 201862
rect 6870 201182 12082 201242
rect 12022 200532 12082 201182
rect 574686 200562 574692 200564
rect 571964 200502 574692 200562
rect 574686 200500 574692 200502
rect 574756 200500 574762 200564
rect 574870 192476 574876 192540
rect 574940 192538 574946 192540
rect 583520 192538 584960 192628
rect 574940 192478 584960 192538
rect 574940 192476 574946 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 6310 188866 6316 188868
rect -960 188806 6316 188866
rect -960 188716 480 188806
rect 6310 188804 6316 188806
rect 6380 188804 6386 188868
rect 6310 186084 6316 186148
rect 6380 186146 6386 186148
rect 574870 186146 574876 186148
rect 6380 186086 12052 186146
rect 571964 186086 574876 186146
rect 6380 186084 6386 186086
rect 574870 186084 574876 186086
rect 574940 186084 574946 186148
rect 574686 179148 574692 179212
rect 574756 179210 574762 179212
rect 583520 179210 584960 179300
rect 574756 179150 584960 179210
rect 574756 179148 574762 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 6310 171668 6316 171732
rect 6380 171730 6386 171732
rect 574686 171730 574692 171732
rect 6380 171670 12052 171730
rect 571964 171670 574692 171730
rect 6380 171668 6386 171670
rect 574686 171668 574692 171670
rect 574756 171668 574762 171732
rect 574870 165820 574876 165884
rect 574940 165882 574946 165884
rect 583520 165882 584960 165972
rect 574940 165822 584960 165882
rect 574940 165820 574946 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 6310 162890 6316 162892
rect -960 162830 6316 162890
rect -960 162740 480 162830
rect 6310 162828 6316 162830
rect 6380 162828 6386 162892
rect 6310 157252 6316 157316
rect 6380 157314 6386 157316
rect 574870 157314 574876 157316
rect 6380 157254 12052 157314
rect 571964 157254 574876 157314
rect 6380 157252 6386 157254
rect 574870 157252 574876 157254
rect 574940 157252 574946 157316
rect 574686 152628 574692 152692
rect 574756 152690 574762 152692
rect 583520 152690 584960 152780
rect 574756 152630 584960 152690
rect 574756 152628 574762 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 6310 149834 6316 149836
rect -960 149774 6316 149834
rect -960 149684 480 149774
rect 6310 149772 6316 149774
rect 6380 149772 6386 149836
rect 4838 142836 4844 142900
rect 4908 142898 4914 142900
rect 574686 142898 574692 142900
rect 4908 142838 12052 142898
rect 571964 142838 574692 142898
rect 4908 142836 4914 142838
rect 574686 142836 574692 142838
rect 574756 142836 574762 142900
rect 574870 139300 574876 139364
rect 574940 139362 574946 139364
rect 583520 139362 584960 139452
rect 574940 139302 584960 139362
rect 574940 139300 574946 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 4838 136778 4844 136780
rect -960 136718 4844 136778
rect -960 136628 480 136718
rect 4838 136716 4844 136718
rect 4908 136716 4914 136780
rect 3366 128420 3372 128484
rect 3436 128482 3442 128484
rect 574870 128482 574876 128484
rect 3436 128422 12052 128482
rect 571964 128422 574876 128482
rect 3436 128420 3442 128422
rect 574870 128420 574876 128422
rect 574940 128420 574946 128484
rect 574686 125972 574692 126036
rect 574756 126034 574762 126036
rect 583520 126034 584960 126124
rect 574756 125974 584960 126034
rect 574756 125972 574762 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 3550 114004 3556 114068
rect 3620 114066 3626 114068
rect 574686 114066 574692 114068
rect 3620 114006 12052 114066
rect 571964 114006 574692 114066
rect 3620 114004 3626 114006
rect 574686 114004 574692 114006
rect 574756 114004 574762 114068
rect 574870 112780 574876 112844
rect 574940 112842 574946 112844
rect 583520 112842 584960 112932
rect 574940 112782 584960 112842
rect 574940 112780 574946 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3366 110666 3372 110668
rect -960 110606 3372 110666
rect -960 110516 480 110606
rect 3366 110604 3372 110606
rect 3436 110604 3442 110668
rect 8886 99588 8892 99652
rect 8956 99650 8962 99652
rect 574870 99650 574876 99652
rect 8956 99590 12052 99650
rect 571964 99590 574876 99650
rect 8956 99588 8962 99590
rect 574870 99588 574876 99590
rect 574940 99588 574946 99652
rect 574686 99452 574692 99516
rect 574756 99514 574762 99516
rect 583520 99514 584960 99604
rect 574756 99454 584960 99514
rect 574756 99452 574762 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3550 97610 3556 97612
rect -960 97550 3556 97610
rect -960 97460 480 97550
rect 3550 97548 3556 97550
rect 3620 97548 3626 97612
rect 574870 86124 574876 86188
rect 574940 86186 574946 86188
rect 583520 86186 584960 86276
rect 574940 86126 584960 86186
rect 574940 86124 574946 86126
rect 583520 86036 584960 86126
rect 8702 85172 8708 85236
rect 8772 85234 8778 85236
rect 574686 85234 574692 85236
rect 8772 85174 12052 85234
rect 571964 85174 574692 85234
rect 8772 85172 8778 85174
rect 574686 85172 574692 85174
rect 574756 85172 574762 85236
rect -960 84690 480 84780
rect 8886 84690 8892 84692
rect -960 84630 8892 84690
rect -960 84540 480 84630
rect 8886 84628 8892 84630
rect 8956 84628 8962 84692
rect 574686 72932 574692 72996
rect 574756 72994 574762 72996
rect 583520 72994 584960 73084
rect 574756 72934 584960 72994
rect 574756 72932 574762 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 8702 71634 8708 71636
rect -960 71574 8708 71634
rect -960 71484 480 71574
rect 8702 71572 8708 71574
rect 8772 71572 8778 71636
rect 8886 70756 8892 70820
rect 8956 70818 8962 70820
rect 574686 70818 574692 70820
rect 8956 70758 12052 70818
rect 571964 70758 574692 70818
rect 8956 70756 8962 70758
rect 574686 70756 574692 70758
rect 574756 70756 574762 70820
rect 574686 59604 574692 59668
rect 574756 59666 574762 59668
rect 583520 59666 584960 59756
rect 574756 59606 584960 59666
rect 574756 59604 574762 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 8886 58578 8892 58580
rect -960 58518 8892 58578
rect -960 58428 480 58518
rect 8886 58516 8892 58518
rect 8956 58516 8962 58580
rect 8886 56340 8892 56404
rect 8956 56402 8962 56404
rect 574686 56402 574692 56404
rect 8956 56342 12052 56402
rect 571964 56342 574692 56402
rect 8956 56340 8962 56342
rect 574686 56340 574692 56342
rect 574756 56340 574762 56404
rect 574686 46276 574692 46340
rect 574756 46338 574762 46340
rect 583520 46338 584960 46428
rect 574756 46278 584960 46338
rect 574756 46276 574762 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 8886 45522 8892 45524
rect -960 45462 8892 45522
rect -960 45372 480 45462
rect 8886 45460 8892 45462
rect 8956 45460 8962 45524
rect 8886 41924 8892 41988
rect 8956 41986 8962 41988
rect 574686 41986 574692 41988
rect 8956 41926 12052 41986
rect 571964 41926 574692 41986
rect 8956 41924 8962 41926
rect 574686 41924 574692 41926
rect 574756 41924 574762 41988
rect 574686 33084 574692 33148
rect 574756 33146 574762 33148
rect 583520 33146 584960 33236
rect 574756 33086 584960 33146
rect 574756 33084 574762 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 8886 32466 8892 32468
rect -960 32406 8892 32466
rect -960 32316 480 32406
rect 8886 32404 8892 32406
rect 8956 32404 8962 32468
rect 6310 27508 6316 27572
rect 6380 27570 6386 27572
rect 575422 27570 575428 27572
rect 6380 27510 12052 27570
rect 571964 27510 575428 27570
rect 6380 27508 6386 27510
rect 575422 27508 575428 27510
rect 575492 27508 575498 27572
rect 575422 19756 575428 19820
rect 575492 19818 575498 19820
rect 583520 19818 584960 19908
rect 575492 19758 584960 19818
rect 575492 19756 575498 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 6310 19410 6316 19412
rect -960 19350 6316 19410
rect -960 19260 480 19350
rect 6310 19348 6316 19350
rect 6380 19348 6386 19412
rect 8886 13092 8892 13156
rect 8956 13154 8962 13156
rect 574686 13154 574692 13156
rect 8956 13094 12052 13154
rect 571964 13094 574692 13154
rect 8956 13092 8962 13094
rect 574686 13092 574692 13094
rect 574756 13092 574762 13156
rect -960 6490 480 6580
rect 574686 6564 574692 6628
rect 574756 6626 574762 6628
rect 583520 6626 584960 6716
rect 574756 6566 584960 6626
rect 574756 6564 574762 6566
rect 8886 6490 8892 6492
rect -960 6430 8892 6490
rect -960 6340 480 6430
rect 8886 6428 8892 6430
rect 8956 6428 8962 6492
rect 583520 6476 584960 6566
rect 47894 3844 47900 3908
rect 47964 3906 47970 3908
rect 59854 3906 59860 3908
rect 47964 3846 59860 3906
rect 47964 3844 47970 3846
rect 59854 3844 59860 3846
rect 59924 3844 59930 3908
rect 558494 3906 558500 3908
rect 553350 3846 558500 3906
rect 383510 3708 383516 3772
rect 383580 3770 383586 3772
rect 389398 3770 389404 3772
rect 383580 3710 389404 3770
rect 383580 3708 383586 3710
rect 389398 3708 389404 3710
rect 389468 3708 389474 3772
rect 533470 3770 533476 3772
rect 526302 3710 533476 3770
rect 526302 3636 526362 3710
rect 533470 3708 533476 3710
rect 533540 3708 533546 3772
rect 462630 3634 462636 3636
rect 452886 3574 462636 3634
rect 397494 3362 397500 3364
rect 392166 3302 397500 3362
rect 34830 3164 34836 3228
rect 34900 3226 34906 3228
rect 34900 3166 45570 3226
rect 34900 3164 34906 3166
rect 35847 2954 35913 2957
rect 17174 2952 35913 2954
rect 17174 2896 35852 2952
rect 35908 2896 35913 2952
rect 17174 2894 35913 2896
rect 45510 2954 45570 3166
rect 364190 3090 364196 3092
rect 55170 3030 66914 3090
rect 52407 2954 52473 2957
rect 55170 2954 55230 3030
rect 66854 2954 66914 3030
rect 363462 3030 364196 3090
rect 68967 2954 69033 2957
rect 45510 2952 52473 2954
rect 45510 2896 52412 2952
rect 52468 2896 52473 2952
rect 45510 2894 52473 2896
rect 17033 2818 17099 2821
rect 17174 2818 17234 2894
rect 35847 2891 35913 2894
rect 52407 2891 52473 2894
rect 53054 2894 55230 2954
rect 58574 2894 64890 2954
rect 66854 2952 69033 2954
rect 66854 2896 68972 2952
rect 69028 2896 69033 2952
rect 66854 2894 69033 2896
rect 17033 2816 17234 2818
rect 17033 2760 17038 2816
rect 17094 2760 17234 2816
rect 17033 2758 17234 2760
rect 23013 2818 23079 2821
rect 41367 2818 41433 2821
rect 23013 2816 41433 2818
rect 23013 2760 23018 2816
rect 23074 2760 41372 2816
rect 41428 2760 41433 2816
rect 23013 2758 41433 2760
rect 17033 2755 17099 2758
rect 23013 2755 23079 2758
rect 41367 2755 41433 2758
rect 41646 2758 52930 2818
rect 40769 2682 40835 2685
rect 41646 2682 41706 2758
rect 47853 2684 47919 2685
rect 47853 2682 47900 2684
rect 40769 2680 41706 2682
rect 40769 2624 40774 2680
rect 40830 2624 41706 2680
rect 40769 2622 41706 2624
rect 47808 2680 47900 2682
rect 47808 2624 47858 2680
rect 47808 2622 47900 2624
rect 40769 2619 40835 2622
rect 47853 2620 47900 2622
rect 47964 2620 47970 2684
rect 47853 2619 47919 2620
rect 34789 2548 34855 2549
rect 34789 2546 34836 2548
rect 34744 2544 34836 2546
rect 34744 2488 34794 2544
rect 34744 2486 34836 2488
rect 34789 2484 34836 2486
rect 34900 2484 34906 2548
rect 52870 2546 52930 2758
rect 53054 2685 53114 2894
rect 57927 2818 57993 2821
rect 53005 2680 53114 2685
rect 53005 2624 53010 2680
rect 53066 2624 53114 2680
rect 53005 2622 53114 2624
rect 53238 2816 57993 2818
rect 53238 2760 57932 2816
rect 57988 2760 57993 2816
rect 53238 2758 57993 2760
rect 53005 2619 53071 2622
rect 53238 2546 53298 2758
rect 57927 2755 57993 2758
rect 58433 2818 58499 2821
rect 58574 2818 58634 2894
rect 58433 2816 58634 2818
rect 58433 2760 58438 2816
rect 58494 2760 58634 2816
rect 58433 2758 58634 2760
rect 58433 2755 58499 2758
rect 59854 2756 59860 2820
rect 59924 2818 59930 2820
rect 64321 2818 64387 2821
rect 59924 2816 64387 2818
rect 59924 2760 64326 2816
rect 64382 2760 64387 2816
rect 59924 2758 64387 2760
rect 64830 2818 64890 2894
rect 68967 2891 69033 2894
rect 74487 2952 74553 2957
rect 74487 2896 74492 2952
rect 74548 2896 74553 2952
rect 74487 2891 74553 2896
rect 353799 2954 353865 2957
rect 360423 2954 360489 2957
rect 363462 2954 363522 3030
rect 364190 3028 364196 3030
rect 364260 3028 364266 3092
rect 377438 3090 377444 3092
rect 372662 3030 377444 3090
rect 353799 2952 356898 2954
rect 353799 2896 353804 2952
rect 353860 2896 356898 2952
rect 353799 2894 356898 2896
rect 353799 2891 353865 2894
rect 74490 2818 74550 2891
rect 356838 2821 356898 2894
rect 357390 2894 360210 2954
rect 64830 2758 74550 2818
rect 76189 2818 76255 2821
rect 91047 2818 91113 2821
rect 76189 2816 91113 2818
rect 76189 2760 76194 2816
rect 76250 2760 91052 2816
rect 91108 2760 91113 2816
rect 76189 2758 91113 2760
rect 59924 2756 59930 2758
rect 64321 2755 64387 2758
rect 76189 2755 76255 2758
rect 91047 2755 91113 2758
rect 91553 2818 91619 2821
rect 105399 2818 105465 2821
rect 91553 2816 105465 2818
rect 91553 2760 91558 2816
rect 91614 2760 105404 2816
rect 105460 2760 105465 2816
rect 91553 2758 105465 2760
rect 91553 2755 91619 2758
rect 105399 2755 105465 2758
rect 117681 2818 117747 2821
rect 129687 2818 129753 2821
rect 117681 2816 129753 2818
rect 117681 2760 117686 2816
rect 117742 2760 129692 2816
rect 129748 2760 129753 2816
rect 117681 2758 129753 2760
rect 117681 2755 117747 2758
rect 129687 2755 129753 2758
rect 147121 2818 147187 2821
rect 157287 2818 157353 2821
rect 147121 2816 157353 2818
rect 147121 2760 147126 2816
rect 147182 2760 157292 2816
rect 157348 2760 157353 2816
rect 147121 2758 157353 2760
rect 147121 2755 147187 2758
rect 157287 2755 157353 2758
rect 186129 2818 186195 2821
rect 193719 2818 193785 2821
rect 186129 2816 193785 2818
rect 186129 2760 186134 2816
rect 186190 2760 193724 2816
rect 193780 2760 193785 2816
rect 186129 2758 193785 2760
rect 186129 2755 186195 2758
rect 193719 2755 193785 2758
rect 344967 2818 345033 2821
rect 346071 2818 346137 2821
rect 349245 2818 349311 2821
rect 344967 2816 345858 2818
rect 344967 2760 344972 2816
rect 345028 2760 345858 2816
rect 344967 2758 345858 2760
rect 344967 2755 345033 2758
rect 109309 2682 109375 2685
rect 121913 2682 121979 2685
rect 109309 2680 121979 2682
rect 109309 2624 109314 2680
rect 109370 2624 121918 2680
rect 121974 2624 121979 2680
rect 109309 2622 121979 2624
rect 109309 2619 109375 2622
rect 121913 2619 121979 2622
rect 150617 2682 150683 2685
rect 160553 2682 160619 2685
rect 150617 2680 160619 2682
rect 150617 2624 150622 2680
rect 150678 2624 160558 2680
rect 160614 2624 160619 2680
rect 150617 2622 160619 2624
rect 150617 2619 150683 2622
rect 160553 2619 160619 2622
rect 218053 2682 218119 2685
rect 223481 2682 223547 2685
rect 218053 2680 223547 2682
rect 218053 2624 218058 2680
rect 218114 2624 223486 2680
rect 223542 2624 223547 2680
rect 218053 2622 223547 2624
rect 345798 2682 345858 2758
rect 346071 2816 349311 2818
rect 346071 2760 346076 2816
rect 346132 2760 349250 2816
rect 349306 2760 349311 2816
rect 346071 2758 349311 2760
rect 346071 2755 346137 2758
rect 349245 2755 349311 2758
rect 350487 2818 350553 2821
rect 352695 2818 352761 2821
rect 356329 2818 356395 2821
rect 350487 2816 352482 2818
rect 350487 2760 350492 2816
rect 350548 2760 352482 2816
rect 350487 2758 352482 2760
rect 350487 2755 350553 2758
rect 347773 2682 347839 2685
rect 345798 2680 347839 2682
rect 345798 2624 347778 2680
rect 347834 2624 347839 2680
rect 345798 2622 347839 2624
rect 352422 2682 352482 2758
rect 352695 2816 356395 2818
rect 352695 2760 352700 2816
rect 352756 2760 356334 2816
rect 356390 2760 356395 2816
rect 352695 2758 356395 2760
rect 356838 2816 356947 2821
rect 356838 2760 356886 2816
rect 356942 2760 356947 2816
rect 356838 2758 356947 2760
rect 352695 2755 352761 2758
rect 356329 2755 356395 2758
rect 356881 2755 356947 2758
rect 357111 2818 357177 2821
rect 357390 2818 357450 2894
rect 359917 2818 359983 2821
rect 357111 2816 357450 2818
rect 357111 2760 357116 2816
rect 357172 2760 357450 2816
rect 357111 2758 357450 2760
rect 357758 2816 359983 2818
rect 357758 2760 359922 2816
rect 359978 2760 359983 2816
rect 357758 2758 359983 2760
rect 360150 2818 360210 2894
rect 360423 2952 363522 2954
rect 360423 2896 360428 2952
rect 360484 2896 363522 2952
rect 360423 2894 363522 2896
rect 363735 2954 363801 2957
rect 363735 2952 368122 2954
rect 363735 2896 363740 2952
rect 363796 2896 368122 2952
rect 363735 2894 368122 2896
rect 360423 2891 360489 2894
rect 363735 2891 363801 2894
rect 361113 2818 361179 2821
rect 360150 2816 361179 2818
rect 360150 2760 361118 2816
rect 361174 2760 361179 2816
rect 360150 2758 361179 2760
rect 357111 2755 357177 2758
rect 353293 2682 353359 2685
rect 352422 2680 353359 2682
rect 352422 2624 353298 2680
rect 353354 2624 353359 2680
rect 352422 2622 353359 2624
rect 218053 2619 218119 2622
rect 223481 2619 223547 2622
rect 347773 2619 347839 2622
rect 353293 2619 353359 2622
rect 356053 2682 356119 2685
rect 357758 2682 357818 2758
rect 359917 2755 359983 2758
rect 361113 2755 361179 2758
rect 361527 2818 361593 2821
rect 364057 2818 364123 2821
rect 361527 2816 364123 2818
rect 361527 2760 361532 2816
rect 361588 2760 364062 2816
rect 364118 2760 364123 2816
rect 361527 2758 364123 2760
rect 361527 2755 361593 2758
rect 364057 2755 364123 2758
rect 364190 2756 364196 2820
rect 364260 2818 364266 2820
rect 364609 2818 364675 2821
rect 364260 2816 364675 2818
rect 364260 2760 364614 2816
rect 364670 2760 364675 2816
rect 364260 2758 364675 2760
rect 364260 2756 364266 2758
rect 364609 2755 364675 2758
rect 364839 2818 364905 2821
rect 368062 2818 368122 2894
rect 368197 2818 368263 2821
rect 364839 2816 367938 2818
rect 364839 2760 364844 2816
rect 364900 2760 367938 2816
rect 364839 2758 367938 2760
rect 368062 2816 368263 2818
rect 368062 2760 368202 2816
rect 368258 2760 368263 2816
rect 368062 2758 368263 2760
rect 364839 2755 364905 2758
rect 356053 2680 357818 2682
rect 356053 2624 356058 2680
rect 356114 2624 357818 2680
rect 356053 2622 357818 2624
rect 367878 2682 367938 2758
rect 368197 2755 368263 2758
rect 369255 2818 369321 2821
rect 371325 2818 371391 2821
rect 369255 2816 371391 2818
rect 369255 2760 369260 2816
rect 369316 2760 371330 2816
rect 371386 2760 371391 2816
rect 369255 2758 371391 2760
rect 369255 2755 369321 2758
rect 371325 2755 371391 2758
rect 371463 2818 371529 2821
rect 372521 2818 372587 2821
rect 372662 2818 372722 3030
rect 377438 3028 377444 3030
rect 377508 3028 377514 3092
rect 383610 3030 387810 3090
rect 373671 2954 373737 2957
rect 382503 2954 382569 2957
rect 383610 2954 383670 3030
rect 373671 2952 378794 2954
rect 373671 2896 373676 2952
rect 373732 2896 378794 2952
rect 373671 2894 378794 2896
rect 373671 2891 373737 2894
rect 376477 2818 376543 2821
rect 378734 2818 378794 2894
rect 382503 2952 383670 2954
rect 382503 2896 382508 2952
rect 382564 2896 383670 2952
rect 382503 2894 383670 2896
rect 383886 2894 387074 2954
rect 382503 2891 382569 2894
rect 378869 2818 378935 2821
rect 371463 2816 372354 2818
rect 371463 2760 371468 2816
rect 371524 2760 372354 2816
rect 371463 2758 372354 2760
rect 371463 2755 371529 2758
rect 369025 2682 369091 2685
rect 367878 2680 369091 2682
rect 367878 2624 369030 2680
rect 369086 2624 369091 2680
rect 367878 2622 369091 2624
rect 372294 2682 372354 2758
rect 372521 2816 372722 2818
rect 372521 2760 372526 2816
rect 372582 2760 372722 2816
rect 372521 2758 372722 2760
rect 372846 2816 376543 2818
rect 372846 2760 376482 2816
rect 376538 2760 376543 2816
rect 372846 2758 376543 2760
rect 372521 2755 372587 2758
rect 372846 2682 372906 2758
rect 376477 2755 376543 2758
rect 376710 2758 378610 2818
rect 378734 2816 378935 2818
rect 378734 2760 378874 2816
rect 378930 2760 378935 2816
rect 378734 2758 378935 2760
rect 372294 2622 372906 2682
rect 374821 2682 374887 2685
rect 376710 2682 376770 2758
rect 374821 2680 376770 2682
rect 374821 2624 374826 2680
rect 374882 2624 376770 2680
rect 374821 2622 376770 2624
rect 378550 2682 378610 2758
rect 378869 2755 378935 2758
rect 379191 2818 379257 2821
rect 381399 2818 381465 2821
rect 383886 2818 383946 2894
rect 384757 2818 384823 2821
rect 379191 2816 381186 2818
rect 379191 2760 379196 2816
rect 379252 2760 381186 2816
rect 379191 2758 381186 2760
rect 379191 2755 379257 2758
rect 379513 2682 379579 2685
rect 378550 2680 379579 2682
rect 378550 2624 379518 2680
rect 379574 2624 379579 2680
rect 378550 2622 379579 2624
rect 381126 2682 381186 2758
rect 381399 2816 383946 2818
rect 381399 2760 381404 2816
rect 381460 2760 383946 2816
rect 381399 2758 383946 2760
rect 384070 2816 384823 2818
rect 384070 2760 384762 2816
rect 384818 2760 384823 2816
rect 384070 2758 384823 2760
rect 381399 2755 381465 2758
rect 384070 2682 384130 2758
rect 384757 2755 384823 2758
rect 384941 2818 385007 2821
rect 387014 2818 387074 2894
rect 387750 2821 387810 3030
rect 391335 2954 391401 2957
rect 392166 2954 392226 3302
rect 397494 3300 397500 3302
rect 397564 3300 397570 3364
rect 405958 3226 405964 3228
rect 401366 3166 405964 3226
rect 391335 2952 392226 2954
rect 391335 2896 391340 2952
rect 391396 2896 392226 2952
rect 391335 2894 392226 2896
rect 392439 2954 392505 2957
rect 399063 2954 399129 2957
rect 401366 2954 401426 3166
rect 405958 3164 405964 3166
rect 406028 3164 406034 3228
rect 402930 3030 408786 3090
rect 392439 2952 398666 2954
rect 392439 2896 392444 2952
rect 392500 2896 398666 2952
rect 392439 2894 398666 2896
rect 391335 2891 391401 2894
rect 392439 2891 392505 2894
rect 387149 2818 387215 2821
rect 384941 2816 386890 2818
rect 384941 2760 384946 2816
rect 385002 2760 386890 2816
rect 384941 2758 386890 2760
rect 387014 2816 387215 2818
rect 387014 2760 387154 2816
rect 387210 2760 387215 2816
rect 387014 2758 387215 2760
rect 387750 2816 387859 2821
rect 387750 2760 387798 2816
rect 387854 2760 387859 2816
rect 387750 2758 387859 2760
rect 384941 2755 385007 2758
rect 381126 2622 384130 2682
rect 386830 2682 386890 2758
rect 387149 2755 387215 2758
rect 387793 2755 387859 2758
rect 388023 2818 388089 2821
rect 393221 2818 393287 2821
rect 388023 2816 393287 2818
rect 388023 2760 388028 2816
rect 388084 2760 393226 2816
rect 393282 2760 393287 2816
rect 388023 2758 393287 2760
rect 388023 2755 388089 2758
rect 393221 2755 393287 2758
rect 393497 2818 393563 2821
rect 395337 2818 395403 2821
rect 393497 2816 395403 2818
rect 393497 2760 393502 2816
rect 393558 2760 395342 2816
rect 395398 2760 395403 2816
rect 393497 2758 395403 2760
rect 393497 2755 393563 2758
rect 395337 2755 395403 2758
rect 396855 2818 396921 2821
rect 396855 2816 398482 2818
rect 396855 2760 396860 2816
rect 396916 2760 398482 2816
rect 396855 2758 398482 2760
rect 396855 2755 396921 2758
rect 390553 2682 390619 2685
rect 397545 2684 397611 2685
rect 386830 2680 390619 2682
rect 386830 2624 390558 2680
rect 390614 2624 390619 2680
rect 386830 2622 390619 2624
rect 356053 2619 356119 2622
rect 369025 2619 369091 2622
rect 374821 2619 374887 2622
rect 379513 2619 379579 2622
rect 390553 2619 390619 2622
rect 397494 2620 397500 2684
rect 397564 2682 397611 2684
rect 397564 2680 397656 2682
rect 397606 2624 397656 2680
rect 397564 2622 397656 2624
rect 397564 2620 397611 2622
rect 397545 2619 397611 2620
rect 52870 2486 53298 2546
rect 72601 2546 72667 2549
rect 87689 2546 87755 2549
rect 72601 2544 87755 2546
rect 72601 2488 72606 2544
rect 72662 2488 87694 2544
rect 87750 2488 87755 2544
rect 72601 2486 87755 2488
rect 34789 2483 34855 2484
rect 72601 2483 72667 2486
rect 87689 2483 87755 2486
rect 105721 2546 105787 2549
rect 118601 2546 118667 2549
rect 105721 2544 118667 2546
rect 105721 2488 105726 2544
rect 105782 2488 118606 2544
rect 118662 2488 118667 2544
rect 105721 2486 118667 2488
rect 105721 2483 105787 2486
rect 118601 2483 118667 2486
rect 149513 2546 149579 2549
rect 159449 2546 159515 2549
rect 149513 2544 159515 2546
rect 149513 2488 149518 2544
rect 149574 2488 159454 2544
rect 159510 2488 159515 2544
rect 149513 2486 159515 2488
rect 149513 2483 149579 2486
rect 159449 2483 159515 2486
rect 162485 2546 162551 2549
rect 171593 2546 171659 2549
rect 377489 2548 377555 2549
rect 383561 2548 383627 2549
rect 389449 2548 389515 2549
rect 162485 2544 171659 2546
rect 162485 2488 162490 2544
rect 162546 2488 171598 2544
rect 171654 2488 171659 2544
rect 162485 2486 171659 2488
rect 162485 2483 162551 2486
rect 171593 2483 171659 2486
rect 377438 2484 377444 2548
rect 377508 2546 377555 2548
rect 383510 2546 383516 2548
rect 377508 2544 377600 2546
rect 377550 2488 377600 2544
rect 377508 2486 377600 2488
rect 383470 2486 383516 2546
rect 383580 2544 383627 2548
rect 383622 2488 383627 2544
rect 377508 2484 377555 2486
rect 383510 2484 383516 2486
rect 383580 2484 383627 2488
rect 389398 2484 389404 2548
rect 389468 2546 389515 2548
rect 398422 2546 398482 2758
rect 398606 2682 398666 2894
rect 399063 2952 401426 2954
rect 399063 2896 399068 2952
rect 399124 2896 401426 2952
rect 399063 2894 401426 2896
rect 402375 2954 402441 2957
rect 402930 2954 402990 3030
rect 402375 2952 402990 2954
rect 402375 2896 402380 2952
rect 402436 2896 402990 2952
rect 402375 2894 402990 2896
rect 403479 2954 403545 2957
rect 403479 2952 408602 2954
rect 403479 2896 403484 2952
rect 403540 2896 408602 2952
rect 403479 2894 408602 2896
rect 399063 2891 399129 2894
rect 402375 2891 402441 2894
rect 403479 2891 403545 2894
rect 403617 2818 403683 2821
rect 406009 2820 406075 2821
rect 398974 2816 403683 2818
rect 398974 2760 403622 2816
rect 403678 2760 403683 2816
rect 398974 2758 403683 2760
rect 398833 2682 398899 2685
rect 398606 2680 398899 2682
rect 398606 2624 398838 2680
rect 398894 2624 398899 2680
rect 398606 2622 398899 2624
rect 398833 2619 398899 2622
rect 398974 2546 399034 2758
rect 403617 2755 403683 2758
rect 405958 2756 405964 2820
rect 406028 2818 406075 2820
rect 406028 2816 406120 2818
rect 406070 2760 406120 2816
rect 406028 2758 406120 2760
rect 406028 2756 406075 2758
rect 406009 2755 406075 2756
rect 408542 2682 408602 2894
rect 408726 2818 408786 3030
rect 408999 2954 409065 2957
rect 421143 2954 421209 2957
rect 452055 2954 452121 2957
rect 452886 2954 452946 3574
rect 462630 3572 462636 3574
rect 462700 3572 462706 3636
rect 517830 3634 517836 3636
rect 509190 3574 517836 3634
rect 463734 3498 463740 3500
rect 455094 3438 463740 3498
rect 408999 2952 414858 2954
rect 408999 2896 409004 2952
rect 409060 2896 414858 2952
rect 408999 2894 414858 2896
rect 408999 2891 409065 2894
rect 409597 2818 409663 2821
rect 408726 2816 409663 2818
rect 408726 2760 409602 2816
rect 409658 2760 409663 2816
rect 408726 2758 409663 2760
rect 409597 2755 409663 2758
rect 410103 2818 410169 2821
rect 414798 2818 414858 2894
rect 421143 2952 429210 2954
rect 421143 2896 421148 2952
rect 421204 2896 429210 2952
rect 421143 2894 429210 2896
rect 421143 2891 421209 2894
rect 416589 2818 416655 2821
rect 417969 2818 418035 2821
rect 410103 2816 414674 2818
rect 410103 2760 410108 2816
rect 410164 2760 414674 2816
rect 410103 2758 414674 2760
rect 414798 2816 416655 2818
rect 414798 2760 416594 2816
rect 416650 2760 416655 2816
rect 414798 2758 416655 2760
rect 410103 2755 410169 2758
rect 410425 2682 410491 2685
rect 408542 2680 410491 2682
rect 408542 2624 410430 2680
rect 410486 2624 410491 2680
rect 408542 2622 410491 2624
rect 414614 2682 414674 2758
rect 416589 2755 416655 2758
rect 416822 2816 418035 2818
rect 416822 2760 417974 2816
rect 418030 2760 418035 2816
rect 416822 2758 418035 2760
rect 416822 2682 416882 2758
rect 417969 2755 418035 2758
rect 423351 2818 423417 2821
rect 423351 2816 429026 2818
rect 423351 2760 423356 2816
rect 423412 2760 429026 2816
rect 423351 2758 429026 2760
rect 423351 2755 423417 2758
rect 414614 2622 416882 2682
rect 410425 2619 410491 2622
rect 389468 2544 389560 2546
rect 389510 2488 389560 2544
rect 389468 2486 389560 2488
rect 398422 2486 399034 2546
rect 428966 2546 429026 2758
rect 429150 2685 429210 2894
rect 452055 2952 452946 2954
rect 452055 2896 452060 2952
rect 452116 2896 452946 2952
rect 452055 2894 452946 2896
rect 453159 2954 453225 2957
rect 455094 2954 455154 3438
rect 463734 3436 463740 3438
rect 463804 3436 463810 3500
rect 458398 3300 458404 3364
rect 458468 3362 458474 3364
rect 467230 3362 467236 3364
rect 458468 3302 467236 3362
rect 458468 3300 458474 3302
rect 467230 3300 467236 3302
rect 467300 3300 467306 3364
rect 470550 3302 471162 3362
rect 466310 3226 466316 3228
rect 455370 3166 466316 3226
rect 455370 2957 455430 3166
rect 466310 3164 466316 3166
rect 466380 3164 466386 3228
rect 470550 3226 470610 3302
rect 466502 3166 470610 3226
rect 466502 3090 466562 3166
rect 463926 3030 466562 3090
rect 467054 3030 470610 3090
rect 453159 2952 455154 2954
rect 453159 2896 453164 2952
rect 453220 2896 455154 2952
rect 453159 2894 455154 2896
rect 455367 2952 455433 2957
rect 455367 2896 455372 2952
rect 455428 2896 455433 2952
rect 452055 2891 452121 2894
rect 453159 2891 453225 2894
rect 455367 2891 455433 2896
rect 456471 2954 456537 2957
rect 458398 2954 458404 2956
rect 456471 2952 458404 2954
rect 456471 2896 456476 2952
rect 456532 2896 458404 2952
rect 456471 2894 458404 2896
rect 456471 2891 456537 2894
rect 458398 2892 458404 2894
rect 458468 2892 458474 2956
rect 458679 2954 458745 2957
rect 459783 2954 459849 2957
rect 463926 2954 463986 3030
rect 458679 2952 459570 2954
rect 458679 2896 458684 2952
rect 458740 2896 459570 2952
rect 458679 2894 459570 2896
rect 458679 2891 458745 2894
rect 432045 2818 432111 2821
rect 429334 2816 432111 2818
rect 429334 2760 432050 2816
rect 432106 2760 432111 2816
rect 429334 2758 432111 2760
rect 459510 2818 459570 2894
rect 459783 2952 463986 2954
rect 459783 2896 459788 2952
rect 459844 2896 463986 2952
rect 459783 2894 463986 2896
rect 464199 2954 464265 2957
rect 467054 2954 467114 3030
rect 464199 2952 467114 2954
rect 464199 2896 464204 2952
rect 464260 2896 467114 2952
rect 464199 2894 467114 2896
rect 459783 2891 459849 2894
rect 464199 2891 464265 2894
rect 459510 2758 463618 2818
rect 429150 2680 429259 2685
rect 429150 2624 429198 2680
rect 429254 2624 429259 2680
rect 429150 2622 429259 2624
rect 429193 2619 429259 2622
rect 429334 2546 429394 2758
rect 432045 2755 432111 2758
rect 441061 2682 441127 2685
rect 450905 2682 450971 2685
rect 462681 2684 462747 2685
rect 441061 2680 450971 2682
rect 441061 2624 441066 2680
rect 441122 2624 450910 2680
rect 450966 2624 450971 2680
rect 441061 2622 450971 2624
rect 441061 2619 441127 2622
rect 450905 2619 450971 2622
rect 462630 2620 462636 2684
rect 462700 2682 462747 2684
rect 463558 2682 463618 2758
rect 463734 2756 463740 2820
rect 463804 2818 463810 2820
rect 463969 2818 464035 2821
rect 469857 2818 469923 2821
rect 463804 2816 464035 2818
rect 463804 2760 463974 2816
rect 464030 2760 464035 2816
rect 463804 2758 464035 2760
rect 463804 2756 463810 2758
rect 463969 2755 464035 2758
rect 464294 2816 469923 2818
rect 464294 2760 469862 2816
rect 469918 2760 469923 2816
rect 464294 2758 469923 2760
rect 470550 2818 470610 3030
rect 471102 2821 471162 3302
rect 498142 3090 498148 3092
rect 489870 3030 498148 3090
rect 471927 2954 471993 2957
rect 485175 2954 485241 2957
rect 489870 2954 489930 3030
rect 498142 3028 498148 3030
rect 498212 3028 498218 3092
rect 471927 2952 483858 2954
rect 471927 2896 471932 2952
rect 471988 2896 483858 2952
rect 471927 2894 483858 2896
rect 471927 2891 471993 2894
rect 470550 2758 470978 2818
rect 464294 2682 464354 2758
rect 469857 2755 469923 2758
rect 462700 2680 462792 2682
rect 462742 2624 462792 2680
rect 462700 2622 462792 2624
rect 463558 2622 464354 2682
rect 470918 2682 470978 2758
rect 471053 2816 471162 2821
rect 471053 2760 471058 2816
rect 471114 2760 471162 2816
rect 471053 2758 471162 2760
rect 471237 2818 471303 2821
rect 482829 2818 482895 2821
rect 471237 2816 482895 2818
rect 471237 2760 471242 2816
rect 471298 2760 482834 2816
rect 482890 2760 482895 2816
rect 471237 2758 482895 2760
rect 483798 2818 483858 2894
rect 485175 2952 489930 2954
rect 485175 2896 485180 2952
rect 485236 2896 489930 2952
rect 485175 2894 489930 2896
rect 495111 2954 495177 2957
rect 508359 2954 508425 2957
rect 509190 2954 509250 3574
rect 517830 3572 517836 3574
rect 517900 3572 517906 3636
rect 526294 3572 526300 3636
rect 526364 3572 526370 3636
rect 545246 3634 545252 3636
rect 530718 3574 545252 3634
rect 516726 3436 516732 3500
rect 516796 3498 516802 3500
rect 516796 3438 530042 3498
rect 516796 3436 516802 3438
rect 517102 3302 527650 3362
rect 514518 3164 514524 3228
rect 514588 3226 514594 3228
rect 517102 3226 517162 3302
rect 514588 3166 517162 3226
rect 517470 3166 524430 3226
rect 514588 3164 514594 3166
rect 495111 2952 508146 2954
rect 495111 2896 495116 2952
rect 495172 2896 508146 2952
rect 495111 2894 508146 2896
rect 485175 2891 485241 2894
rect 495111 2891 495177 2894
rect 483933 2818 483999 2821
rect 483798 2816 483999 2818
rect 483798 2760 483938 2816
rect 483994 2760 483999 2816
rect 483798 2758 483999 2760
rect 471053 2755 471119 2758
rect 471237 2755 471303 2758
rect 482829 2755 482895 2758
rect 483933 2755 483999 2758
rect 491799 2818 491865 2821
rect 505369 2818 505435 2821
rect 491799 2816 505435 2818
rect 491799 2760 491804 2816
rect 491860 2760 505374 2816
rect 505430 2760 505435 2816
rect 491799 2758 505435 2760
rect 508086 2818 508146 2894
rect 508359 2952 509250 2954
rect 508359 2896 508364 2952
rect 508420 2896 509250 2952
rect 508359 2894 509250 2896
rect 511671 2954 511737 2957
rect 514983 2954 515049 2957
rect 516726 2954 516732 2956
rect 511671 2952 514770 2954
rect 511671 2896 511676 2952
rect 511732 2896 514770 2952
rect 511671 2894 514770 2896
rect 508359 2891 508425 2894
rect 511671 2891 511737 2894
rect 508865 2818 508931 2821
rect 508086 2816 508931 2818
rect 508086 2760 508870 2816
rect 508926 2760 508931 2816
rect 508086 2758 508931 2760
rect 491799 2755 491865 2758
rect 505369 2755 505435 2758
rect 508865 2755 508931 2758
rect 509463 2818 509529 2821
rect 512775 2818 512841 2821
rect 514518 2818 514524 2820
rect 509463 2816 512562 2818
rect 509463 2760 509468 2816
rect 509524 2760 512562 2816
rect 509463 2758 512562 2760
rect 509463 2755 509529 2758
rect 475377 2682 475443 2685
rect 470918 2680 475443 2682
rect 470918 2624 475382 2680
rect 475438 2624 475443 2680
rect 470918 2622 475443 2624
rect 512502 2682 512562 2758
rect 512775 2816 514524 2818
rect 512775 2760 512780 2816
rect 512836 2760 514524 2816
rect 512775 2758 514524 2760
rect 512775 2755 512841 2758
rect 514518 2756 514524 2758
rect 514588 2756 514594 2820
rect 514710 2818 514770 2894
rect 514983 2952 516732 2954
rect 514983 2896 514988 2952
rect 515044 2896 516732 2952
rect 514983 2894 516732 2896
rect 514983 2891 515049 2894
rect 516726 2892 516732 2894
rect 516796 2892 516802 2956
rect 517470 2954 517530 3166
rect 517830 3028 517836 3092
rect 517900 3090 517906 3092
rect 522982 3090 522988 3092
rect 517900 3030 522988 3090
rect 517900 3028 517906 3030
rect 522982 3028 522988 3030
rect 523052 3028 523058 3092
rect 524370 3090 524430 3166
rect 527590 3092 527650 3302
rect 529982 3228 530042 3438
rect 529974 3164 529980 3228
rect 530044 3164 530050 3228
rect 526478 3090 526484 3092
rect 524370 3030 526484 3090
rect 526478 3028 526484 3030
rect 526548 3028 526554 3092
rect 527582 3028 527588 3092
rect 527652 3028 527658 3092
rect 517102 2894 517530 2954
rect 518295 2954 518361 2957
rect 524919 2954 524985 2957
rect 526294 2954 526300 2956
rect 518295 2952 524430 2954
rect 518295 2896 518300 2952
rect 518356 2896 524430 2952
rect 518295 2894 524430 2896
rect 517102 2818 517162 2894
rect 518295 2891 518361 2894
rect 524229 2818 524295 2821
rect 514710 2758 517162 2818
rect 517286 2816 524295 2818
rect 517286 2760 524234 2816
rect 524290 2760 524295 2816
rect 517286 2758 524295 2760
rect 524370 2818 524430 2894
rect 524919 2952 526300 2954
rect 524919 2896 524924 2952
rect 524980 2896 526300 2952
rect 524919 2894 526300 2896
rect 524919 2891 524985 2894
rect 526294 2892 526300 2894
rect 526364 2892 526370 2956
rect 529335 2954 529401 2957
rect 530718 2954 530778 3574
rect 545246 3572 545252 3574
rect 545316 3572 545322 3636
rect 547638 3498 547644 3500
rect 534950 3438 543750 3498
rect 533340 3030 534090 3090
rect 529335 2952 530778 2954
rect 529335 2896 529340 2952
rect 529396 2896 530778 2952
rect 529335 2894 530778 2896
rect 531543 2954 531609 2957
rect 533340 2954 533400 3030
rect 531543 2952 533400 2954
rect 531543 2896 531548 2952
rect 531604 2896 533400 2952
rect 531543 2894 533400 2896
rect 529335 2891 529401 2894
rect 531543 2891 531609 2894
rect 533470 2892 533476 2956
rect 533540 2892 533546 2956
rect 534030 2954 534090 3030
rect 534950 2954 535010 3438
rect 543690 3362 543750 3438
rect 545438 3438 547644 3498
rect 545438 3362 545498 3438
rect 547638 3436 547644 3438
rect 547708 3436 547714 3500
rect 552422 3362 552428 3364
rect 543690 3302 545498 3362
rect 547462 3302 552428 3362
rect 547462 3226 547522 3302
rect 552422 3300 552428 3302
rect 552492 3300 552498 3364
rect 553350 3226 553410 3846
rect 558494 3844 558500 3846
rect 558564 3844 558570 3908
rect 538170 3166 547522 3226
rect 547830 3166 553410 3226
rect 534030 2894 535010 2954
rect 535959 2954 536025 2957
rect 538170 2954 538230 3166
rect 535959 2952 538230 2954
rect 535959 2896 535964 2952
rect 536020 2896 538230 2952
rect 535959 2894 538230 2896
rect 541479 2954 541545 2957
rect 547830 2954 547890 3166
rect 557490 3030 562058 3090
rect 541479 2952 547890 2954
rect 541479 2896 541484 2952
rect 541540 2896 547890 2952
rect 541479 2894 547890 2896
rect 548103 2954 548169 2957
rect 557490 2954 557550 3030
rect 548103 2952 557550 2954
rect 548103 2896 548108 2952
rect 548164 2896 557550 2952
rect 548103 2894 557550 2896
rect 533286 2818 533292 2820
rect 524370 2758 533292 2818
rect 517286 2682 517346 2758
rect 524229 2755 524295 2758
rect 533286 2756 533292 2758
rect 533356 2756 533362 2820
rect 533478 2818 533538 2892
rect 535959 2891 536025 2894
rect 541479 2891 541545 2894
rect 548103 2891 548169 2894
rect 540789 2818 540855 2821
rect 533478 2816 540855 2818
rect 533478 2760 540794 2816
rect 540850 2760 540855 2816
rect 533478 2758 540855 2760
rect 540789 2755 540855 2758
rect 542583 2818 542649 2821
rect 558545 2820 558611 2821
rect 542583 2816 558378 2818
rect 542583 2760 542588 2816
rect 542644 2760 558378 2816
rect 542583 2758 558378 2760
rect 542583 2755 542649 2758
rect 526529 2684 526595 2685
rect 527633 2684 527699 2685
rect 530025 2684 530091 2685
rect 533337 2684 533403 2685
rect 552473 2684 552539 2685
rect 512502 2622 517346 2682
rect 462700 2620 462747 2622
rect 462681 2619 462747 2620
rect 475377 2619 475443 2622
rect 526478 2620 526484 2684
rect 526548 2682 526595 2684
rect 526548 2680 526640 2682
rect 526590 2624 526640 2680
rect 526548 2622 526640 2624
rect 526548 2620 526595 2622
rect 527582 2620 527588 2684
rect 527652 2682 527699 2684
rect 527652 2680 527744 2682
rect 527694 2624 527744 2680
rect 527652 2622 527744 2624
rect 527652 2620 527699 2622
rect 529974 2620 529980 2684
rect 530044 2682 530091 2684
rect 530044 2680 530136 2682
rect 530086 2624 530136 2680
rect 530044 2622 530136 2624
rect 530044 2620 530091 2622
rect 533286 2620 533292 2684
rect 533356 2682 533403 2684
rect 533356 2680 533448 2682
rect 533398 2624 533448 2680
rect 533356 2622 533448 2624
rect 533356 2620 533403 2622
rect 552422 2620 552428 2684
rect 552492 2682 552539 2684
rect 552492 2680 552584 2682
rect 552534 2624 552584 2680
rect 552492 2622 552584 2624
rect 552492 2620 552539 2622
rect 526529 2619 526595 2620
rect 527633 2619 527699 2620
rect 530025 2619 530091 2620
rect 533337 2619 533403 2620
rect 552473 2619 552539 2620
rect 428966 2486 429394 2546
rect 430021 2546 430087 2549
rect 439129 2546 439195 2549
rect 430021 2544 439195 2546
rect 430021 2488 430026 2544
rect 430082 2488 439134 2544
rect 439190 2488 439195 2544
rect 430021 2486 439195 2488
rect 389468 2484 389515 2486
rect 377489 2483 377555 2484
rect 383561 2483 383627 2484
rect 389449 2483 389515 2484
rect 430021 2483 430087 2486
rect 439129 2483 439195 2486
rect 442165 2546 442231 2549
rect 452101 2546 452167 2549
rect 466269 2548 466335 2549
rect 467281 2548 467347 2549
rect 498193 2548 498259 2549
rect 523033 2548 523099 2549
rect 545297 2548 545363 2549
rect 466269 2546 466316 2548
rect 442165 2544 452167 2546
rect 442165 2488 442170 2544
rect 442226 2488 452106 2544
rect 452162 2488 452167 2544
rect 442165 2486 452167 2488
rect 466224 2544 466316 2546
rect 466224 2488 466274 2544
rect 466224 2486 466316 2488
rect 442165 2483 442231 2486
rect 452101 2483 452167 2486
rect 466269 2484 466316 2486
rect 466380 2484 466386 2548
rect 467230 2484 467236 2548
rect 467300 2546 467347 2548
rect 467300 2544 467392 2546
rect 467342 2488 467392 2544
rect 467300 2486 467392 2488
rect 467300 2484 467347 2486
rect 498142 2484 498148 2548
rect 498212 2546 498259 2548
rect 498212 2544 498304 2546
rect 498254 2488 498304 2544
rect 498212 2486 498304 2488
rect 498212 2484 498259 2486
rect 522982 2484 522988 2548
rect 523052 2546 523099 2548
rect 523052 2544 523144 2546
rect 523094 2488 523144 2544
rect 523052 2486 523144 2488
rect 523052 2484 523099 2486
rect 545246 2484 545252 2548
rect 545316 2546 545363 2548
rect 545316 2544 545408 2546
rect 545358 2488 545408 2544
rect 545316 2486 545408 2488
rect 545316 2484 545363 2486
rect 547638 2484 547644 2548
rect 547708 2546 547714 2548
rect 547873 2546 547939 2549
rect 547708 2544 547939 2546
rect 547708 2488 547878 2544
rect 547934 2488 547939 2544
rect 547708 2486 547939 2488
rect 558318 2546 558378 2758
rect 558494 2756 558500 2820
rect 558564 2818 558611 2820
rect 561998 2818 562058 3030
rect 565629 2818 565695 2821
rect 558564 2816 558656 2818
rect 558606 2760 558656 2816
rect 558564 2758 558656 2760
rect 561998 2816 565695 2818
rect 561998 2760 565634 2816
rect 565690 2760 565695 2816
rect 561998 2758 565695 2760
rect 558564 2756 558611 2758
rect 558545 2755 558611 2756
rect 565629 2755 565695 2758
rect 559281 2546 559347 2549
rect 558318 2544 559347 2546
rect 558318 2488 559286 2544
rect 559342 2488 559347 2544
rect 558318 2486 559347 2488
rect 547708 2484 547714 2486
rect 466269 2483 466335 2484
rect 467281 2483 467347 2484
rect 498193 2483 498259 2484
rect 523033 2483 523099 2484
rect 545297 2483 545363 2484
rect 547873 2483 547939 2486
rect 559281 2483 559347 2486
rect 69105 2410 69171 2413
rect 84377 2410 84443 2413
rect 69105 2408 84443 2410
rect 69105 2352 69110 2408
rect 69166 2352 84382 2408
rect 84438 2352 84443 2408
rect 69105 2350 84443 2352
rect 69105 2347 69171 2350
rect 84377 2347 84443 2350
rect 102225 2410 102291 2413
rect 115289 2410 115355 2413
rect 102225 2408 115355 2410
rect 102225 2352 102230 2408
rect 102286 2352 115294 2408
rect 115350 2352 115355 2408
rect 102225 2350 115355 2352
rect 102225 2347 102291 2350
rect 115289 2347 115355 2350
rect 143533 2410 143599 2413
rect 153929 2410 153995 2413
rect 143533 2408 153995 2410
rect 143533 2352 143538 2408
rect 143594 2352 153934 2408
rect 153990 2352 153995 2408
rect 143533 2350 153995 2352
rect 143533 2347 143599 2350
rect 153929 2347 153995 2350
rect 156597 2410 156663 2413
rect 166073 2410 166139 2413
rect 156597 2408 166139 2410
rect 156597 2352 156602 2408
rect 156658 2352 166078 2408
rect 166134 2352 166139 2408
rect 156597 2350 166139 2352
rect 156597 2347 156663 2350
rect 166073 2347 166139 2350
rect 216857 2410 216923 2413
rect 222377 2410 222443 2413
rect 216857 2408 222443 2410
rect 216857 2352 216862 2408
rect 216918 2352 222382 2408
rect 222438 2352 222443 2408
rect 216857 2350 222443 2352
rect 216857 2347 216923 2350
rect 222377 2347 222443 2350
rect 228725 2410 228791 2413
rect 233417 2410 233483 2413
rect 228725 2408 233483 2410
rect 228725 2352 228730 2408
rect 228786 2352 233422 2408
rect 233478 2352 233483 2408
rect 228725 2350 233483 2352
rect 228725 2347 228791 2350
rect 233417 2347 233483 2350
rect 246389 2410 246455 2413
rect 249977 2410 250043 2413
rect 246389 2408 250043 2410
rect 246389 2352 246394 2408
rect 246450 2352 249982 2408
rect 250038 2352 250043 2408
rect 246389 2350 250043 2352
rect 246389 2347 246455 2350
rect 249977 2347 250043 2350
rect 433241 2410 433307 2413
rect 442625 2410 442691 2413
rect 433241 2408 442691 2410
rect 433241 2352 433246 2408
rect 433302 2352 442630 2408
rect 442686 2352 442691 2408
rect 433241 2350 442691 2352
rect 433241 2347 433307 2350
rect 442625 2347 442691 2350
rect 443269 2410 443335 2413
rect 453297 2410 453363 2413
rect 443269 2408 453363 2410
rect 443269 2352 443274 2408
rect 443330 2352 453302 2408
rect 453358 2352 453363 2408
rect 443269 2350 453363 2352
rect 443269 2347 443335 2350
rect 453297 2347 453363 2350
rect 66989 2274 67055 2277
rect 82169 2274 82235 2277
rect 66989 2272 82235 2274
rect 66989 2216 66994 2272
rect 67050 2216 82174 2272
rect 82230 2216 82235 2272
rect 66989 2214 82235 2216
rect 66989 2211 67055 2214
rect 82169 2211 82235 2214
rect 99741 2274 99807 2277
rect 113081 2274 113147 2277
rect 99741 2272 113147 2274
rect 99741 2216 99746 2272
rect 99802 2216 113086 2272
rect 113142 2216 113147 2272
rect 99741 2214 113147 2216
rect 99741 2211 99807 2214
rect 113081 2211 113147 2214
rect 141233 2274 141299 2277
rect 151721 2274 151787 2277
rect 141233 2272 151787 2274
rect 141233 2216 141238 2272
rect 141294 2216 151726 2272
rect 151782 2216 151787 2272
rect 141233 2214 151787 2216
rect 141233 2211 141299 2214
rect 151721 2211 151787 2214
rect 155401 2274 155467 2277
rect 164969 2274 165035 2277
rect 155401 2272 165035 2274
rect 155401 2216 155406 2272
rect 155462 2216 164974 2272
rect 165030 2216 165035 2272
rect 155401 2214 165035 2216
rect 155401 2211 155467 2214
rect 164969 2211 165035 2214
rect 209773 2274 209839 2277
rect 215753 2274 215819 2277
rect 209773 2272 215819 2274
rect 209773 2216 209778 2272
rect 209834 2216 215758 2272
rect 215814 2216 215819 2272
rect 209773 2214 215819 2216
rect 209773 2211 209839 2214
rect 215753 2211 215819 2214
rect 219249 2274 219315 2277
rect 224585 2274 224651 2277
rect 219249 2272 224651 2274
rect 219249 2216 219254 2272
rect 219310 2216 224590 2272
rect 224646 2216 224651 2272
rect 219249 2214 224651 2216
rect 219249 2211 219315 2214
rect 224585 2211 224651 2214
rect 435541 2274 435607 2277
rect 445017 2274 445083 2277
rect 435541 2272 445083 2274
rect 435541 2216 435546 2272
rect 435602 2216 445022 2272
rect 445078 2216 445083 2272
rect 435541 2214 445083 2216
rect 435541 2211 435607 2214
rect 445017 2211 445083 2214
rect 445477 2274 445543 2277
rect 455689 2274 455755 2277
rect 445477 2272 455755 2274
rect 445477 2216 445482 2272
rect 445538 2216 455694 2272
rect 455750 2216 455755 2272
rect 445477 2214 455755 2216
rect 445477 2211 445543 2214
rect 455689 2211 455755 2214
rect 463141 2274 463207 2277
rect 474549 2274 474615 2277
rect 463141 2272 474615 2274
rect 463141 2216 463146 2272
rect 463202 2216 474554 2272
rect 474610 2216 474615 2272
rect 463141 2214 474615 2216
rect 463141 2211 463207 2214
rect 474549 2211 474615 2214
rect 65517 2138 65583 2141
rect 81065 2138 81131 2141
rect 65517 2136 81131 2138
rect 65517 2080 65522 2136
rect 65578 2080 81070 2136
rect 81126 2080 81131 2136
rect 65517 2078 81131 2080
rect 65517 2075 65583 2078
rect 81065 2075 81131 2078
rect 101029 2138 101095 2141
rect 114185 2138 114251 2141
rect 101029 2136 114251 2138
rect 101029 2080 101034 2136
rect 101090 2080 114190 2136
rect 114246 2080 114251 2136
rect 101029 2078 114251 2080
rect 101029 2075 101095 2078
rect 114185 2075 114251 2078
rect 115197 2138 115263 2141
rect 127433 2138 127499 2141
rect 115197 2136 127499 2138
rect 115197 2080 115202 2136
rect 115258 2080 127438 2136
rect 127494 2080 127499 2136
rect 115197 2078 127499 2080
rect 115197 2075 115263 2078
rect 127433 2075 127499 2078
rect 142429 2138 142495 2141
rect 152825 2138 152891 2141
rect 142429 2136 152891 2138
rect 142429 2080 142434 2136
rect 142490 2080 152830 2136
rect 152886 2080 152891 2136
rect 142429 2078 152891 2080
rect 142429 2075 142495 2078
rect 152825 2075 152891 2078
rect 154205 2138 154271 2141
rect 163865 2138 163931 2141
rect 154205 2136 163931 2138
rect 154205 2080 154210 2136
rect 154266 2080 163870 2136
rect 163926 2080 163931 2136
rect 154205 2078 163931 2080
rect 154205 2075 154271 2078
rect 163865 2075 163931 2078
rect 207381 2138 207447 2141
rect 213545 2138 213611 2141
rect 207381 2136 213611 2138
rect 207381 2080 207386 2136
rect 207442 2080 213550 2136
rect 213606 2080 213611 2136
rect 207381 2078 213611 2080
rect 207381 2075 207447 2078
rect 213545 2075 213611 2078
rect 223941 2138 224007 2141
rect 229001 2138 229067 2141
rect 223941 2136 229067 2138
rect 223941 2080 223946 2136
rect 224002 2080 229006 2136
rect 229062 2080 229067 2136
rect 223941 2078 229067 2080
rect 223941 2075 224007 2078
rect 229001 2075 229067 2078
rect 229829 2138 229895 2141
rect 234521 2138 234587 2141
rect 229829 2136 234587 2138
rect 229829 2080 229834 2136
rect 229890 2080 234526 2136
rect 234582 2080 234587 2136
rect 229829 2078 234587 2080
rect 229829 2075 229895 2078
rect 234521 2075 234587 2078
rect 239305 2138 239371 2141
rect 243353 2138 243419 2141
rect 239305 2136 243419 2138
rect 239305 2080 239310 2136
rect 239366 2080 243358 2136
rect 243414 2080 243419 2136
rect 239305 2078 243419 2080
rect 239305 2075 239371 2078
rect 243353 2075 243419 2078
rect 424501 2138 424567 2141
rect 433241 2138 433307 2141
rect 424501 2136 433307 2138
rect 424501 2080 424506 2136
rect 424562 2080 433246 2136
rect 433302 2080 433307 2136
rect 424501 2078 433307 2080
rect 424501 2075 424567 2078
rect 433241 2075 433307 2078
rect 436645 2138 436711 2141
rect 446213 2138 446279 2141
rect 436645 2136 446279 2138
rect 436645 2080 436650 2136
rect 436706 2080 446218 2136
rect 446274 2080 446279 2136
rect 436645 2078 446279 2080
rect 436645 2075 436711 2078
rect 446213 2075 446279 2078
rect 446581 2138 446647 2141
rect 456885 2138 456951 2141
rect 446581 2136 456951 2138
rect 446581 2080 446586 2136
rect 446642 2080 456890 2136
rect 456946 2080 456951 2136
rect 446581 2078 456951 2080
rect 446581 2075 446647 2078
rect 456885 2075 456951 2078
rect 468661 2138 468727 2141
rect 480529 2138 480595 2141
rect 468661 2136 480595 2138
rect 468661 2080 468666 2136
rect 468722 2080 480534 2136
rect 480590 2080 480595 2136
rect 468661 2078 480595 2080
rect 468661 2075 468727 2078
rect 480529 2075 480595 2078
rect 59629 2002 59695 2005
rect 75545 2002 75611 2005
rect 59629 2000 75611 2002
rect 59629 1944 59634 2000
rect 59690 1944 75550 2000
rect 75606 1944 75611 2000
rect 59629 1942 75611 1944
rect 59629 1939 59695 1942
rect 75545 1939 75611 1942
rect 93945 2002 94011 2005
rect 107561 2002 107627 2005
rect 93945 2000 107627 2002
rect 93945 1944 93950 2000
rect 94006 1944 107566 2000
rect 107622 1944 107627 2000
rect 93945 1942 107627 1944
rect 93945 1939 94011 1942
rect 107561 1939 107627 1942
rect 108113 2002 108179 2005
rect 120809 2002 120875 2005
rect 108113 2000 120875 2002
rect 108113 1944 108118 2000
rect 108174 1944 120814 2000
rect 120870 1944 120875 2000
rect 108113 1942 120875 1944
rect 108113 1939 108179 1942
rect 120809 1939 120875 1942
rect 135253 2002 135319 2005
rect 146201 2002 146267 2005
rect 135253 2000 146267 2002
rect 135253 1944 135258 2000
rect 135314 1944 146206 2000
rect 146262 1944 146267 2000
rect 135253 1942 146267 1944
rect 135253 1939 135319 1942
rect 146201 1939 146267 1942
rect 148317 2002 148383 2005
rect 158345 2002 158411 2005
rect 148317 2000 158411 2002
rect 148317 1944 148322 2000
rect 148378 1944 158350 2000
rect 158406 1944 158411 2000
rect 148317 1942 158411 1944
rect 148317 1939 148383 1942
rect 158345 1939 158411 1942
rect 161289 2002 161355 2005
rect 170489 2002 170555 2005
rect 161289 2000 170555 2002
rect 161289 1944 161294 2000
rect 161350 1944 170494 2000
rect 170550 1944 170555 2000
rect 161289 1942 170555 1944
rect 161289 1939 161355 1942
rect 170489 1939 170555 1942
rect 180241 2002 180307 2005
rect 188153 2002 188219 2005
rect 180241 2000 188219 2002
rect 180241 1944 180246 2000
rect 180302 1944 188158 2000
rect 188214 1944 188219 2000
rect 180241 1942 188219 1944
rect 180241 1939 180307 1942
rect 188153 1939 188219 1942
rect 189717 2002 189783 2005
rect 196985 2002 197051 2005
rect 189717 2000 197051 2002
rect 189717 1944 189722 2000
rect 189778 1944 196990 2000
rect 197046 1944 197051 2000
rect 189717 1942 197051 1944
rect 189717 1939 189783 1942
rect 196985 1939 197051 1942
rect 208577 2002 208643 2005
rect 214649 2002 214715 2005
rect 208577 2000 214715 2002
rect 208577 1944 208582 2000
rect 208638 1944 214654 2000
rect 214710 1944 214715 2000
rect 208577 1942 214715 1944
rect 208577 1939 208643 1942
rect 214649 1939 214715 1942
rect 220445 2002 220511 2005
rect 225689 2002 225755 2005
rect 220445 2000 225755 2002
rect 220445 1944 220450 2000
rect 220506 1944 225694 2000
rect 225750 1944 225755 2000
rect 220445 1942 225755 1944
rect 220445 1939 220511 1942
rect 225689 1939 225755 1942
rect 227529 2002 227595 2005
rect 232313 2002 232379 2005
rect 227529 2000 232379 2002
rect 227529 1944 227534 2000
rect 227590 1944 232318 2000
rect 232374 1944 232379 2000
rect 227529 1942 232379 1944
rect 227529 1939 227595 1942
rect 232313 1939 232379 1942
rect 238109 2002 238175 2005
rect 242249 2002 242315 2005
rect 238109 2000 242315 2002
rect 238109 1944 238114 2000
rect 238170 1944 242254 2000
rect 242310 1944 242315 2000
rect 238109 1942 242315 1944
rect 238109 1939 238175 1942
rect 242249 1939 242315 1942
rect 248781 2002 248847 2005
rect 252185 2002 252251 2005
rect 248781 2000 252251 2002
rect 248781 1944 248786 2000
rect 248842 1944 252190 2000
rect 252246 1944 252251 2000
rect 248781 1942 252251 1944
rect 248781 1939 248847 1942
rect 252185 1939 252251 1942
rect 401317 2002 401383 2005
rect 408401 2002 408467 2005
rect 401317 2000 408467 2002
rect 401317 1944 401322 2000
rect 401378 1944 408406 2000
rect 408462 1944 408467 2000
rect 401317 1942 408467 1944
rect 401317 1939 401383 1942
rect 408401 1939 408467 1942
rect 418981 2002 419047 2005
rect 427261 2002 427327 2005
rect 418981 2000 427327 2002
rect 418981 1944 418986 2000
rect 419042 1944 427266 2000
rect 427322 1944 427327 2000
rect 418981 1942 427327 1944
rect 418981 1939 419047 1942
rect 427261 1939 427327 1942
rect 427721 2002 427787 2005
rect 436737 2002 436803 2005
rect 427721 2000 436803 2002
rect 427721 1944 427726 2000
rect 427782 1944 436742 2000
rect 436798 1944 436803 2000
rect 427721 1942 436803 1944
rect 427721 1939 427787 1942
rect 436737 1939 436803 1942
rect 437749 2002 437815 2005
rect 447409 2002 447475 2005
rect 437749 2000 447475 2002
rect 437749 1944 437754 2000
rect 437810 1944 447414 2000
rect 447470 1944 447475 2000
rect 437749 1942 447475 1944
rect 437749 1939 437815 1942
rect 447409 1939 447475 1942
rect 448789 2002 448855 2005
rect 459185 2002 459251 2005
rect 448789 2000 459251 2002
rect 448789 1944 448794 2000
rect 448850 1944 459190 2000
rect 459246 1944 459251 2000
rect 448789 1942 459251 1944
rect 448789 1939 448855 1942
rect 459185 1939 459251 1942
rect 469765 2002 469831 2005
rect 481725 2002 481791 2005
rect 469765 2000 481791 2002
rect 469765 1944 469770 2000
rect 469826 1944 481730 2000
rect 481786 1944 481791 2000
rect 469765 1942 481791 1944
rect 469765 1939 469831 1942
rect 481725 1939 481791 1942
rect 528277 2002 528343 2005
rect 544377 2002 544443 2005
rect 528277 2000 544443 2002
rect 528277 1944 528282 2000
rect 528338 1944 544382 2000
rect 544438 1944 544443 2000
rect 528277 1942 544443 1944
rect 528277 1939 528343 1942
rect 544377 1939 544443 1942
rect 111609 1866 111675 1869
rect 124121 1866 124187 1869
rect 111609 1864 124187 1866
rect 111609 1808 111614 1864
rect 111670 1808 124126 1864
rect 124182 1808 124187 1864
rect 111609 1806 124187 1808
rect 111609 1803 111675 1806
rect 124121 1803 124187 1806
rect 151813 1866 151879 1869
rect 161657 1866 161723 1869
rect 151813 1864 161723 1866
rect 151813 1808 151818 1864
rect 151874 1808 161662 1864
rect 161718 1808 161723 1864
rect 151813 1806 161723 1808
rect 151813 1803 151879 1806
rect 161657 1803 161723 1806
rect 212165 1866 212231 1869
rect 217961 1866 218027 1869
rect 212165 1864 218027 1866
rect 212165 1808 212170 1864
rect 212226 1808 217966 1864
rect 218022 1808 218027 1864
rect 212165 1806 218027 1808
rect 212165 1803 212231 1806
rect 217961 1803 218027 1806
rect 221549 1866 221615 1869
rect 226793 1866 226859 1869
rect 221549 1864 226859 1866
rect 221549 1808 221554 1864
rect 221610 1808 226798 1864
rect 226854 1808 226859 1864
rect 221549 1806 226859 1808
rect 221549 1803 221615 1806
rect 226793 1803 226859 1806
rect 233417 1866 233483 1869
rect 237833 1866 237899 1869
rect 233417 1864 237899 1866
rect 233417 1808 233422 1864
rect 233478 1808 237838 1864
rect 237894 1808 237899 1864
rect 233417 1806 237899 1808
rect 233417 1803 233483 1806
rect 237833 1803 237899 1806
rect 241697 1866 241763 1869
rect 245561 1866 245627 1869
rect 241697 1864 245627 1866
rect 241697 1808 241702 1864
rect 241758 1808 245566 1864
rect 245622 1808 245627 1864
rect 241697 1806 245627 1808
rect 241697 1803 241763 1806
rect 245561 1803 245627 1806
rect 247585 1866 247651 1869
rect 251081 1866 251147 1869
rect 247585 1864 251147 1866
rect 247585 1808 247590 1864
rect 247646 1808 251086 1864
rect 251142 1808 251147 1864
rect 247585 1806 251147 1808
rect 247585 1803 247651 1806
rect 251081 1803 251147 1806
rect 439957 1866 440023 1869
rect 449801 1866 449867 1869
rect 439957 1864 449867 1866
rect 439957 1808 439962 1864
rect 440018 1808 449806 1864
rect 449862 1808 449867 1864
rect 439957 1806 449867 1808
rect 439957 1803 440023 1806
rect 449801 1803 449867 1806
rect 112805 1730 112871 1733
rect 125225 1730 125291 1733
rect 112805 1728 125291 1730
rect 112805 1672 112810 1728
rect 112866 1672 125230 1728
rect 125286 1672 125291 1728
rect 112805 1670 125291 1672
rect 112805 1667 112871 1670
rect 125225 1667 125291 1670
rect 157793 1730 157859 1733
rect 167177 1730 167243 1733
rect 157793 1728 167243 1730
rect 157793 1672 157798 1728
rect 157854 1672 167182 1728
rect 167238 1672 167243 1728
rect 157793 1670 167243 1672
rect 157793 1667 157859 1670
rect 167177 1667 167243 1670
rect 200481 1730 200547 1733
rect 206921 1730 206987 1733
rect 200481 1728 206987 1730
rect 200481 1672 200486 1728
rect 200542 1672 206926 1728
rect 206982 1672 206987 1728
rect 200481 1670 206987 1672
rect 200481 1667 200547 1670
rect 206921 1667 206987 1670
rect 213361 1730 213427 1733
rect 219065 1730 219131 1733
rect 213361 1728 219131 1730
rect 213361 1672 213366 1728
rect 213422 1672 219070 1728
rect 219126 1672 219131 1728
rect 213361 1670 219131 1672
rect 213361 1667 213427 1670
rect 219065 1667 219131 1670
rect 222745 1730 222811 1733
rect 227897 1730 227963 1733
rect 222745 1728 227963 1730
rect 222745 1672 222750 1728
rect 222806 1672 227902 1728
rect 227958 1672 227963 1728
rect 222745 1670 227963 1672
rect 222745 1667 222811 1670
rect 227897 1667 227963 1670
rect 234613 1730 234679 1733
rect 238937 1730 239003 1733
rect 234613 1728 239003 1730
rect 234613 1672 234618 1728
rect 234674 1672 238942 1728
rect 238998 1672 239003 1728
rect 234613 1670 239003 1672
rect 234613 1667 234679 1670
rect 238937 1667 239003 1670
rect 242893 1730 242959 1733
rect 246665 1730 246731 1733
rect 242893 1728 246731 1730
rect 242893 1672 242898 1728
rect 242954 1672 246670 1728
rect 246726 1672 246731 1728
rect 242893 1670 246731 1672
rect 242893 1667 242959 1670
rect 246665 1667 246731 1670
rect 251173 1730 251239 1733
rect 254393 1730 254459 1733
rect 251173 1728 254459 1730
rect 251173 1672 251178 1728
rect 251234 1672 254398 1728
rect 254454 1672 254459 1728
rect 251173 1670 254459 1672
rect 251173 1667 251239 1670
rect 254393 1667 254459 1670
rect 254669 1730 254735 1733
rect 257705 1730 257771 1733
rect 254669 1728 257771 1730
rect 254669 1672 254674 1728
rect 254730 1672 257710 1728
rect 257766 1672 257771 1728
rect 254669 1670 257771 1672
rect 254669 1667 254735 1670
rect 257705 1667 257771 1670
rect 258257 1730 258323 1733
rect 261017 1730 261083 1733
rect 258257 1728 261083 1730
rect 258257 1672 258262 1728
rect 258318 1672 261022 1728
rect 261078 1672 261083 1728
rect 258257 1670 261083 1672
rect 258257 1667 258323 1670
rect 261017 1667 261083 1670
rect 261753 1730 261819 1733
rect 264329 1730 264395 1733
rect 261753 1728 264395 1730
rect 261753 1672 261758 1728
rect 261814 1672 264334 1728
rect 264390 1672 264395 1728
rect 261753 1670 264395 1672
rect 261753 1667 261819 1670
rect 264329 1667 264395 1670
rect 434437 1730 434503 1733
rect 443821 1730 443887 1733
rect 434437 1728 443887 1730
rect 434437 1672 434442 1728
rect 434498 1672 443826 1728
rect 443882 1672 443887 1728
rect 434437 1670 443887 1672
rect 434437 1667 434503 1670
rect 443821 1667 443887 1670
rect 206185 1594 206251 1597
rect 212441 1594 212507 1597
rect 206185 1592 212507 1594
rect 206185 1536 206190 1592
rect 206246 1536 212446 1592
rect 212502 1536 212507 1592
rect 206185 1534 212507 1536
rect 206185 1531 206251 1534
rect 212441 1531 212507 1534
rect 215661 1594 215727 1597
rect 221273 1594 221339 1597
rect 215661 1592 221339 1594
rect 215661 1536 215666 1592
rect 215722 1536 221278 1592
rect 221334 1536 221339 1592
rect 215661 1534 221339 1536
rect 215661 1531 215727 1534
rect 221273 1531 221339 1534
rect 226333 1594 226399 1597
rect 231209 1594 231275 1597
rect 226333 1592 231275 1594
rect 226333 1536 226338 1592
rect 226394 1536 231214 1592
rect 231270 1536 231275 1592
rect 226333 1534 231275 1536
rect 226333 1531 226399 1534
rect 231209 1531 231275 1534
rect 232221 1594 232287 1597
rect 236729 1594 236795 1597
rect 232221 1592 236795 1594
rect 232221 1536 232226 1592
rect 232282 1536 236734 1592
rect 236790 1536 236795 1592
rect 232221 1534 236795 1536
rect 232221 1531 232287 1534
rect 236729 1531 236795 1534
rect 237005 1594 237071 1597
rect 241145 1594 241211 1597
rect 237005 1592 241211 1594
rect 237005 1536 237010 1592
rect 237066 1536 241150 1592
rect 241206 1536 241211 1592
rect 237005 1534 241211 1536
rect 237005 1531 237071 1534
rect 241145 1531 241211 1534
rect 244089 1594 244155 1597
rect 247769 1594 247835 1597
rect 244089 1592 247835 1594
rect 244089 1536 244094 1592
rect 244150 1536 247774 1592
rect 247830 1536 247835 1592
rect 244089 1534 247835 1536
rect 244089 1531 244155 1534
rect 247769 1531 247835 1534
rect 249977 1594 250043 1597
rect 253289 1594 253355 1597
rect 249977 1592 253355 1594
rect 249977 1536 249982 1592
rect 250038 1536 253294 1592
rect 253350 1536 253355 1592
rect 249977 1534 253355 1536
rect 249977 1531 250043 1534
rect 253289 1531 253355 1534
rect 253473 1594 253539 1597
rect 256601 1594 256667 1597
rect 253473 1592 256667 1594
rect 253473 1536 253478 1592
rect 253534 1536 256606 1592
rect 256662 1536 256667 1592
rect 253473 1534 256667 1536
rect 253473 1531 253539 1534
rect 256601 1531 256667 1534
rect 257061 1594 257127 1597
rect 259913 1594 259979 1597
rect 257061 1592 259979 1594
rect 257061 1536 257066 1592
rect 257122 1536 259918 1592
rect 259974 1536 259979 1592
rect 257061 1534 259979 1536
rect 257061 1531 257127 1534
rect 259913 1531 259979 1534
rect 260649 1594 260715 1597
rect 263225 1594 263291 1597
rect 260649 1592 263291 1594
rect 260649 1536 260654 1592
rect 260710 1536 263230 1592
rect 263286 1536 263291 1592
rect 260649 1534 263291 1536
rect 260649 1531 260715 1534
rect 263225 1531 263291 1534
rect 264145 1594 264211 1597
rect 266537 1594 266603 1597
rect 264145 1592 266603 1594
rect 264145 1536 264150 1592
rect 264206 1536 266542 1592
rect 266598 1536 266603 1592
rect 264145 1534 266603 1536
rect 264145 1531 264211 1534
rect 266537 1531 266603 1534
rect 270033 1594 270099 1597
rect 272057 1594 272123 1597
rect 270033 1592 272123 1594
rect 270033 1536 270038 1592
rect 270094 1536 272062 1592
rect 272118 1536 272123 1592
rect 270033 1534 272123 1536
rect 270033 1531 270099 1534
rect 272057 1531 272123 1534
rect 201493 1458 201559 1461
rect 208025 1458 208091 1461
rect 201493 1456 208091 1458
rect 201493 1400 201498 1456
rect 201554 1400 208030 1456
rect 208086 1400 208091 1456
rect 201493 1398 208091 1400
rect 201493 1395 201559 1398
rect 208025 1395 208091 1398
rect 214465 1458 214531 1461
rect 220169 1458 220235 1461
rect 214465 1456 220235 1458
rect 214465 1400 214470 1456
rect 214526 1400 220174 1456
rect 220230 1400 220235 1456
rect 214465 1398 220235 1400
rect 214465 1395 214531 1398
rect 220169 1395 220235 1398
rect 225137 1458 225203 1461
rect 230105 1458 230171 1461
rect 225137 1456 230171 1458
rect 225137 1400 225142 1456
rect 225198 1400 230110 1456
rect 230166 1400 230171 1456
rect 225137 1398 230171 1400
rect 225137 1395 225203 1398
rect 230105 1395 230171 1398
rect 231025 1458 231091 1461
rect 235625 1458 235691 1461
rect 231025 1456 235691 1458
rect 231025 1400 231030 1456
rect 231086 1400 235630 1456
rect 235686 1400 235691 1456
rect 231025 1398 235691 1400
rect 231025 1395 231091 1398
rect 235625 1395 235691 1398
rect 235809 1458 235875 1461
rect 240041 1458 240107 1461
rect 235809 1456 240107 1458
rect 235809 1400 235814 1456
rect 235870 1400 240046 1456
rect 240102 1400 240107 1456
rect 235809 1398 240107 1400
rect 235809 1395 235875 1398
rect 240041 1395 240107 1398
rect 240501 1458 240567 1461
rect 244457 1458 244523 1461
rect 240501 1456 244523 1458
rect 240501 1400 240506 1456
rect 240562 1400 244462 1456
rect 244518 1400 244523 1456
rect 240501 1398 244523 1400
rect 240501 1395 240567 1398
rect 244457 1395 244523 1398
rect 245193 1458 245259 1461
rect 248873 1458 248939 1461
rect 245193 1456 248939 1458
rect 245193 1400 245198 1456
rect 245254 1400 248878 1456
rect 248934 1400 248939 1456
rect 245193 1398 248939 1400
rect 245193 1395 245259 1398
rect 248873 1395 248939 1398
rect 252369 1458 252435 1461
rect 255497 1458 255563 1461
rect 252369 1456 255563 1458
rect 252369 1400 252374 1456
rect 252430 1400 255502 1456
rect 255558 1400 255563 1456
rect 252369 1398 255563 1400
rect 252369 1395 252435 1398
rect 255497 1395 255563 1398
rect 255865 1458 255931 1461
rect 258809 1458 258875 1461
rect 255865 1456 258875 1458
rect 255865 1400 255870 1456
rect 255926 1400 258814 1456
rect 258870 1400 258875 1456
rect 255865 1398 258875 1400
rect 255865 1395 255931 1398
rect 258809 1395 258875 1398
rect 262949 1458 263015 1461
rect 265433 1458 265499 1461
rect 262949 1456 265499 1458
rect 262949 1400 262954 1456
rect 263010 1400 265438 1456
rect 265494 1400 265499 1456
rect 262949 1398 265499 1400
rect 262949 1395 263015 1398
rect 265433 1395 265499 1398
rect 268837 1458 268903 1461
rect 270953 1458 271019 1461
rect 268837 1456 271019 1458
rect 268837 1400 268842 1456
rect 268898 1400 270958 1456
rect 271014 1400 271019 1456
rect 268837 1398 271019 1400
rect 268837 1395 268903 1398
rect 270953 1395 271019 1398
rect 164877 1322 164943 1325
rect 173801 1322 173867 1325
rect 164877 1320 173867 1322
rect 164877 1264 164882 1320
rect 164938 1264 173806 1320
rect 173862 1264 173867 1320
rect 164877 1262 173867 1264
rect 164877 1259 164943 1262
rect 173801 1259 173867 1262
rect 174261 1322 174327 1325
rect 182633 1322 182699 1325
rect 174261 1320 182699 1322
rect 174261 1264 174266 1320
rect 174322 1264 182638 1320
rect 182694 1264 182699 1320
rect 174261 1262 182699 1264
rect 174261 1259 174327 1262
rect 182633 1259 182699 1262
rect 184933 1322 184999 1325
rect 192569 1322 192635 1325
rect 184933 1320 192635 1322
rect 184933 1264 184938 1320
rect 184994 1264 192574 1320
rect 192630 1264 192635 1320
rect 184933 1262 192635 1264
rect 184933 1259 184999 1262
rect 192569 1259 192635 1262
rect 195605 1322 195671 1325
rect 202505 1322 202571 1325
rect 195605 1320 202571 1322
rect 195605 1264 195610 1320
rect 195666 1264 202510 1320
rect 202566 1264 202571 1320
rect 195605 1262 202571 1264
rect 195605 1259 195671 1262
rect 202505 1259 202571 1262
rect 205081 1322 205147 1325
rect 211337 1322 211403 1325
rect 205081 1320 211403 1322
rect 205081 1264 205086 1320
rect 205142 1264 211342 1320
rect 211398 1264 211403 1320
rect 205081 1262 211403 1264
rect 205081 1259 205147 1262
rect 211337 1259 211403 1262
rect 259453 1322 259519 1325
rect 262121 1322 262187 1325
rect 259453 1320 262187 1322
rect 259453 1264 259458 1320
rect 259514 1264 262126 1320
rect 262182 1264 262187 1320
rect 259453 1262 262187 1264
rect 259453 1259 259519 1262
rect 262121 1259 262187 1262
rect 267733 1322 267799 1325
rect 269849 1322 269915 1325
rect 267733 1320 269915 1322
rect 267733 1264 267738 1320
rect 267794 1264 269854 1320
rect 269910 1264 269915 1320
rect 267733 1262 269915 1264
rect 267733 1259 267799 1262
rect 269849 1259 269915 1262
rect 271229 1322 271295 1325
rect 273161 1322 273227 1325
rect 271229 1320 273227 1322
rect 271229 1264 271234 1320
rect 271290 1264 273166 1320
rect 273222 1264 273227 1320
rect 271229 1262 273227 1264
rect 271229 1259 271295 1262
rect 273161 1259 273227 1262
rect 273621 1322 273687 1325
rect 275369 1322 275435 1325
rect 273621 1320 275435 1322
rect 273621 1264 273626 1320
rect 273682 1264 275374 1320
rect 275430 1264 275435 1320
rect 273621 1262 275435 1264
rect 273621 1259 273687 1262
rect 275369 1259 275435 1262
rect 276013 1322 276079 1325
rect 277577 1322 277643 1325
rect 276013 1320 277643 1322
rect 276013 1264 276018 1320
rect 276074 1264 277582 1320
rect 277638 1264 277643 1320
rect 276013 1262 277643 1264
rect 276013 1259 276079 1262
rect 277577 1259 277643 1262
rect 279509 1322 279575 1325
rect 280889 1322 280955 1325
rect 279509 1320 280955 1322
rect 279509 1264 279514 1320
rect 279570 1264 280894 1320
rect 280950 1264 280955 1320
rect 279509 1262 280955 1264
rect 279509 1259 279575 1262
rect 280889 1259 280955 1262
rect 281901 1322 281967 1325
rect 283189 1322 283255 1325
rect 281901 1320 283255 1322
rect 281901 1264 281906 1320
rect 281962 1264 283194 1320
rect 283250 1264 283255 1320
rect 281901 1262 283255 1264
rect 281901 1259 281967 1262
rect 283189 1259 283255 1262
rect 285397 1322 285463 1325
rect 286409 1322 286475 1325
rect 285397 1320 286475 1322
rect 285397 1264 285402 1320
rect 285458 1264 286414 1320
rect 286470 1264 286475 1320
rect 285397 1262 286475 1264
rect 285397 1259 285463 1262
rect 286409 1259 286475 1262
rect 286593 1322 286659 1325
rect 287513 1322 287579 1325
rect 286593 1320 287579 1322
rect 286593 1264 286598 1320
rect 286654 1264 287518 1320
rect 287574 1264 287579 1320
rect 286593 1262 287579 1264
rect 286593 1259 286659 1262
rect 287513 1259 287579 1262
rect 287789 1322 287855 1325
rect 288617 1322 288683 1325
rect 287789 1320 288683 1322
rect 287789 1264 287794 1320
rect 287850 1264 288622 1320
rect 288678 1264 288683 1320
rect 287789 1262 288683 1264
rect 287789 1259 287855 1262
rect 288617 1259 288683 1262
rect 312997 1322 313063 1325
rect 313825 1322 313891 1325
rect 312997 1320 313891 1322
rect 312997 1264 313002 1320
rect 313058 1264 313830 1320
rect 313886 1264 313891 1320
rect 312997 1262 313891 1264
rect 312997 1259 313063 1262
rect 313825 1259 313891 1262
rect 314101 1322 314167 1325
rect 315021 1322 315087 1325
rect 314101 1320 315087 1322
rect 314101 1264 314106 1320
rect 314162 1264 315026 1320
rect 315082 1264 315087 1320
rect 314101 1262 315087 1264
rect 314101 1259 314167 1262
rect 315021 1259 315087 1262
rect 315205 1322 315271 1325
rect 316217 1322 316283 1325
rect 315205 1320 316283 1322
rect 315205 1264 315210 1320
rect 315266 1264 316222 1320
rect 316278 1264 316283 1320
rect 315205 1262 316283 1264
rect 315205 1259 315271 1262
rect 316217 1259 316283 1262
rect 317413 1322 317479 1325
rect 318517 1322 318583 1325
rect 317413 1320 318583 1322
rect 317413 1264 317418 1320
rect 317474 1264 318522 1320
rect 318578 1264 318583 1320
rect 317413 1262 318583 1264
rect 317413 1259 317479 1262
rect 318517 1259 318583 1262
rect 319621 1322 319687 1325
rect 320909 1322 320975 1325
rect 319621 1320 320975 1322
rect 319621 1264 319626 1320
rect 319682 1264 320914 1320
rect 320970 1264 320975 1320
rect 319621 1262 320975 1264
rect 319621 1259 319687 1262
rect 320909 1259 320975 1262
rect 322841 1322 322907 1325
rect 324405 1322 324471 1325
rect 322841 1320 324471 1322
rect 322841 1264 322846 1320
rect 322902 1264 324410 1320
rect 324466 1264 324471 1320
rect 322841 1262 324471 1264
rect 322841 1259 322907 1262
rect 324405 1259 324471 1262
rect 325141 1322 325207 1325
rect 326797 1322 326863 1325
rect 325141 1320 326863 1322
rect 325141 1264 325146 1320
rect 325202 1264 326802 1320
rect 326858 1264 326863 1320
rect 325141 1262 326863 1264
rect 325141 1259 325207 1262
rect 326797 1259 326863 1262
rect 327349 1322 327415 1325
rect 329189 1322 329255 1325
rect 327349 1320 329255 1322
rect 327349 1264 327354 1320
rect 327410 1264 329194 1320
rect 329250 1264 329255 1320
rect 327349 1262 329255 1264
rect 327349 1259 327415 1262
rect 329189 1259 329255 1262
rect 329557 1322 329623 1325
rect 331581 1322 331647 1325
rect 329557 1320 331647 1322
rect 329557 1264 329562 1320
rect 329618 1264 331586 1320
rect 331642 1264 331647 1320
rect 329557 1262 331647 1264
rect 329557 1259 329623 1262
rect 331581 1259 331647 1262
rect 335077 1322 335143 1325
rect 337469 1322 337535 1325
rect 335077 1320 337535 1322
rect 335077 1264 335082 1320
rect 335138 1264 337474 1320
rect 337530 1264 337535 1320
rect 335077 1262 337535 1264
rect 335077 1259 335143 1262
rect 337469 1259 337535 1262
rect 338389 1322 338455 1325
rect 340965 1322 341031 1325
rect 338389 1320 341031 1322
rect 338389 1264 338394 1320
rect 338450 1264 340970 1320
rect 341026 1264 341031 1320
rect 338389 1262 341031 1264
rect 338389 1259 338455 1262
rect 340965 1259 341031 1262
rect 341701 1322 341767 1325
rect 344553 1322 344619 1325
rect 341701 1320 344619 1322
rect 341701 1264 341706 1320
rect 341762 1264 344558 1320
rect 344614 1264 344619 1320
rect 341701 1262 344619 1264
rect 341701 1259 341767 1262
rect 344553 1259 344619 1262
rect 347221 1322 347287 1325
rect 350441 1322 350507 1325
rect 347221 1320 350507 1322
rect 347221 1264 347226 1320
rect 347282 1264 350446 1320
rect 350502 1264 350507 1320
rect 347221 1262 350507 1264
rect 347221 1259 347287 1262
rect 350441 1259 350507 1262
rect 354949 1322 355015 1325
rect 358721 1322 358787 1325
rect 354949 1320 358787 1322
rect 354949 1264 354954 1320
rect 355010 1264 358726 1320
rect 358782 1264 358787 1320
rect 354949 1262 358787 1264
rect 354949 1259 355015 1262
rect 358721 1259 358787 1262
rect 398005 1322 398071 1325
rect 404813 1322 404879 1325
rect 398005 1320 404879 1322
rect 398005 1264 398010 1320
rect 398066 1264 404818 1320
rect 404874 1264 404879 1320
rect 398005 1262 404879 1264
rect 398005 1259 398071 1262
rect 404813 1259 404879 1262
rect 406837 1322 406903 1325
rect 414289 1322 414355 1325
rect 406837 1320 414355 1322
rect 406837 1264 406842 1320
rect 406898 1264 414294 1320
rect 414350 1264 414355 1320
rect 406837 1262 414355 1264
rect 406837 1259 406903 1262
rect 414289 1259 414355 1262
rect 415669 1322 415735 1325
rect 423765 1322 423831 1325
rect 415669 1320 423831 1322
rect 415669 1264 415674 1320
rect 415730 1264 423770 1320
rect 423826 1264 423831 1320
rect 415669 1262 423831 1264
rect 415669 1259 415735 1262
rect 423765 1259 423831 1262
rect 425605 1322 425671 1325
rect 434437 1322 434503 1325
rect 425605 1320 434503 1322
rect 425605 1264 425610 1320
rect 425666 1264 434442 1320
rect 434498 1264 434503 1320
rect 425605 1262 434503 1264
rect 425605 1259 425671 1262
rect 434437 1259 434503 1262
rect 171961 1186 172027 1189
rect 180425 1186 180491 1189
rect 171961 1184 180491 1186
rect 171961 1128 171966 1184
rect 172022 1128 180430 1184
rect 180486 1128 180491 1184
rect 171961 1126 180491 1128
rect 171961 1123 172027 1126
rect 180425 1123 180491 1126
rect 183737 1186 183803 1189
rect 191465 1186 191531 1189
rect 183737 1184 191531 1186
rect 183737 1128 183742 1184
rect 183798 1128 191470 1184
rect 191526 1128 191531 1184
rect 183737 1126 191531 1128
rect 183737 1123 183803 1126
rect 191465 1123 191531 1126
rect 194409 1186 194475 1189
rect 201401 1186 201467 1189
rect 194409 1184 201467 1186
rect 194409 1128 194414 1184
rect 194470 1128 201406 1184
rect 201462 1128 201467 1184
rect 194409 1126 201467 1128
rect 194409 1123 194475 1126
rect 201401 1123 201467 1126
rect 203885 1186 203951 1189
rect 210233 1186 210299 1189
rect 203885 1184 210299 1186
rect 203885 1128 203890 1184
rect 203946 1128 210238 1184
rect 210294 1128 210299 1184
rect 203885 1126 210299 1128
rect 203885 1123 203951 1126
rect 210233 1123 210299 1126
rect 210969 1186 211035 1189
rect 216949 1186 217015 1189
rect 210969 1184 217015 1186
rect 210969 1128 210974 1184
rect 211030 1128 216954 1184
rect 217010 1128 217015 1184
rect 210969 1126 217015 1128
rect 210969 1123 211035 1126
rect 216949 1123 217015 1126
rect 266537 1186 266603 1189
rect 268745 1186 268811 1189
rect 266537 1184 268811 1186
rect 266537 1128 266542 1184
rect 266598 1128 268750 1184
rect 268806 1128 268811 1184
rect 266537 1126 268811 1128
rect 266537 1123 266603 1126
rect 268745 1123 268811 1126
rect 272425 1186 272491 1189
rect 274265 1186 274331 1189
rect 272425 1184 274331 1186
rect 272425 1128 272430 1184
rect 272486 1128 274270 1184
rect 274326 1128 274331 1184
rect 272425 1126 274331 1128
rect 272425 1123 272491 1126
rect 274265 1123 274331 1126
rect 274817 1186 274883 1189
rect 276473 1186 276539 1189
rect 274817 1184 276539 1186
rect 274817 1128 274822 1184
rect 274878 1128 276478 1184
rect 276534 1128 276539 1184
rect 274817 1126 276539 1128
rect 274817 1123 274883 1126
rect 276473 1123 276539 1126
rect 277117 1186 277183 1189
rect 278681 1186 278747 1189
rect 277117 1184 278747 1186
rect 277117 1128 277122 1184
rect 277178 1128 278686 1184
rect 278742 1128 278747 1184
rect 277117 1126 278747 1128
rect 277117 1123 277183 1126
rect 278681 1123 278747 1126
rect 280705 1186 280771 1189
rect 281993 1186 282059 1189
rect 280705 1184 282059 1186
rect 280705 1128 280710 1184
rect 280766 1128 281998 1184
rect 282054 1128 282059 1184
rect 280705 1126 282059 1128
rect 280705 1123 280771 1126
rect 281993 1123 282059 1126
rect 318425 1186 318491 1189
rect 319713 1186 319779 1189
rect 318425 1184 319779 1186
rect 318425 1128 318430 1184
rect 318486 1128 319718 1184
rect 319774 1128 319779 1184
rect 318425 1126 319779 1128
rect 318425 1123 318491 1126
rect 319713 1123 319779 1126
rect 320725 1186 320791 1189
rect 322105 1186 322171 1189
rect 320725 1184 322171 1186
rect 320725 1128 320730 1184
rect 320786 1128 322110 1184
rect 322166 1128 322171 1184
rect 320725 1126 322171 1128
rect 320725 1123 320791 1126
rect 322105 1123 322171 1126
rect 324037 1186 324103 1189
rect 325601 1186 325667 1189
rect 324037 1184 325667 1186
rect 324037 1128 324042 1184
rect 324098 1128 325606 1184
rect 325662 1128 325667 1184
rect 324037 1126 325667 1128
rect 324037 1123 324103 1126
rect 325601 1123 325667 1126
rect 326245 1186 326311 1189
rect 327993 1186 328059 1189
rect 326245 1184 328059 1186
rect 326245 1128 326250 1184
rect 326306 1128 327998 1184
rect 328054 1128 328059 1184
rect 326245 1126 328059 1128
rect 326245 1123 326311 1126
rect 327993 1123 328059 1126
rect 328361 1186 328427 1189
rect 330385 1186 330451 1189
rect 328361 1184 330451 1186
rect 328361 1128 328366 1184
rect 328422 1128 330390 1184
rect 330446 1128 330451 1184
rect 328361 1126 330451 1128
rect 328361 1123 328427 1126
rect 330385 1123 330451 1126
rect 330661 1186 330727 1189
rect 332685 1186 332751 1189
rect 330661 1184 332751 1186
rect 330661 1128 330666 1184
rect 330722 1128 332690 1184
rect 332746 1128 332751 1184
rect 330661 1126 332751 1128
rect 330661 1123 330727 1126
rect 332685 1123 332751 1126
rect 332869 1186 332935 1189
rect 335077 1186 335143 1189
rect 332869 1184 335143 1186
rect 332869 1128 332874 1184
rect 332930 1128 335082 1184
rect 335138 1128 335143 1184
rect 332869 1126 335143 1128
rect 332869 1123 332935 1126
rect 335077 1123 335143 1126
rect 336181 1186 336247 1189
rect 338665 1186 338731 1189
rect 336181 1184 338731 1186
rect 336181 1128 336186 1184
rect 336242 1128 338670 1184
rect 338726 1128 338731 1184
rect 336181 1126 338731 1128
rect 336181 1123 336247 1126
rect 338665 1123 338731 1126
rect 339401 1186 339467 1189
rect 342161 1186 342227 1189
rect 339401 1184 342227 1186
rect 339401 1128 339406 1184
rect 339462 1128 342166 1184
rect 342222 1128 342227 1184
rect 339401 1126 342227 1128
rect 339401 1123 339467 1126
rect 342161 1123 342227 1126
rect 342805 1186 342871 1189
rect 345749 1186 345815 1189
rect 342805 1184 345815 1186
rect 342805 1128 342810 1184
rect 342866 1128 345754 1184
rect 345810 1128 345815 1184
rect 342805 1126 345815 1128
rect 342805 1123 342871 1126
rect 345749 1123 345815 1126
rect 348325 1186 348391 1189
rect 351637 1186 351703 1189
rect 348325 1184 351703 1186
rect 348325 1128 348330 1184
rect 348386 1128 351642 1184
rect 351698 1128 351703 1184
rect 348325 1126 351703 1128
rect 348325 1123 348391 1126
rect 351637 1123 351703 1126
rect 416681 1186 416747 1189
rect 424961 1186 425027 1189
rect 416681 1184 425027 1186
rect 416681 1128 416686 1184
rect 416742 1128 424966 1184
rect 425022 1128 425027 1184
rect 416681 1126 425027 1128
rect 416681 1123 416747 1126
rect 424961 1123 425027 1126
rect 432229 1186 432295 1189
rect 441521 1186 441587 1189
rect 432229 1184 441587 1186
rect 432229 1128 432234 1184
rect 432290 1128 441526 1184
rect 441582 1128 441587 1184
rect 432229 1126 441587 1128
rect 432229 1123 432295 1126
rect 441521 1123 441587 1126
rect 6453 1050 6519 1053
rect 10961 1050 11027 1053
rect 6453 1048 11027 1050
rect 6453 992 6458 1048
rect 6514 992 10966 1048
rect 11022 992 11027 1048
rect 6453 990 11027 992
rect 6453 987 6519 990
rect 10961 987 11027 990
rect 12341 1050 12407 1053
rect 19241 1050 19307 1053
rect 12341 1048 19307 1050
rect 12341 992 12346 1048
rect 12402 992 19246 1048
rect 19302 992 19307 1048
rect 12341 990 19307 992
rect 12341 987 12407 990
rect 19241 987 19307 990
rect 21817 1050 21883 1053
rect 23841 1050 23907 1053
rect 21817 1048 23907 1050
rect 21817 992 21822 1048
rect 21878 992 23846 1048
rect 23902 992 23907 1048
rect 21817 990 23907 992
rect 21817 987 21883 990
rect 23841 987 23907 990
rect 132769 1050 132835 1053
rect 141785 1050 141851 1053
rect 132769 1048 141851 1050
rect 132769 992 132774 1048
rect 132830 992 141790 1048
rect 141846 992 141851 1048
rect 132769 990 141851 992
rect 132769 987 132835 990
rect 141785 987 141851 990
rect 168373 1050 168439 1053
rect 177113 1050 177179 1053
rect 168373 1048 177179 1050
rect 168373 992 168378 1048
rect 168434 992 177118 1048
rect 177174 992 177179 1048
rect 168373 990 177179 992
rect 168373 987 168439 990
rect 177113 987 177179 990
rect 177849 1050 177915 1053
rect 185945 1050 186011 1053
rect 177849 1048 186011 1050
rect 177849 992 177854 1048
rect 177910 992 185950 1048
rect 186006 992 186011 1048
rect 177849 990 186011 992
rect 177849 987 177915 990
rect 185945 987 186011 990
rect 193213 1050 193279 1053
rect 200297 1050 200363 1053
rect 193213 1048 200363 1050
rect 193213 992 193218 1048
rect 193274 992 200302 1048
rect 200358 992 200363 1048
rect 193213 990 200363 992
rect 193213 987 193279 990
rect 200297 987 200363 990
rect 202689 1050 202755 1053
rect 209129 1050 209195 1053
rect 202689 1048 209195 1050
rect 202689 992 202694 1048
rect 202750 992 209134 1048
rect 209190 992 209195 1048
rect 202689 990 209195 992
rect 202689 987 202755 990
rect 209129 987 209195 990
rect 265341 1050 265407 1053
rect 267641 1050 267707 1053
rect 265341 1048 267707 1050
rect 265341 992 265346 1048
rect 265402 992 267646 1048
rect 267702 992 267707 1048
rect 265341 990 267707 992
rect 265341 987 265407 990
rect 267641 987 267707 990
rect 278313 1050 278379 1053
rect 279785 1050 279851 1053
rect 278313 1048 279851 1050
rect 278313 992 278318 1048
rect 278374 992 279790 1048
rect 279846 992 279851 1048
rect 278313 990 279851 992
rect 278313 987 278379 990
rect 279785 987 279851 990
rect 321829 1050 321895 1053
rect 323301 1050 323367 1053
rect 321829 1048 323367 1050
rect 321829 992 321834 1048
rect 321890 992 323306 1048
rect 323362 992 323367 1048
rect 321829 990 323367 992
rect 321829 987 321895 990
rect 323301 987 323367 990
rect 333881 1050 333947 1053
rect 336273 1050 336339 1053
rect 333881 1048 336339 1050
rect 333881 992 333886 1048
rect 333942 992 336278 1048
rect 336334 992 336339 1048
rect 333881 990 336339 992
rect 333881 987 333947 990
rect 336273 987 336339 990
rect 337285 1050 337351 1053
rect 339861 1050 339927 1053
rect 337285 1048 339927 1050
rect 337285 992 337290 1048
rect 337346 992 339866 1048
rect 339922 992 339927 1048
rect 337285 990 339927 992
rect 337285 987 337351 990
rect 339861 987 339927 990
rect 340597 1050 340663 1053
rect 343357 1050 343423 1053
rect 340597 1048 343423 1050
rect 340597 992 340602 1048
rect 340658 992 343362 1048
rect 343418 992 343423 1048
rect 340597 990 343423 992
rect 340597 987 340663 990
rect 343357 987 343423 990
rect 343909 1050 343975 1053
rect 346945 1050 347011 1053
rect 343909 1048 347011 1050
rect 343909 992 343914 1048
rect 343970 992 346950 1048
rect 347006 992 347011 1048
rect 343909 990 347011 992
rect 343909 987 343975 990
rect 346945 987 347011 990
rect 349429 1050 349495 1053
rect 352833 1050 352899 1053
rect 349429 1048 352899 1050
rect 349429 992 349434 1048
rect 349490 992 352838 1048
rect 352894 992 352899 1048
rect 349429 990 352899 992
rect 349429 987 349495 990
rect 352833 987 352899 990
rect 413461 1050 413527 1053
rect 421373 1050 421439 1053
rect 413461 1048 421439 1050
rect 413461 992 413466 1048
rect 413522 992 421378 1048
rect 421434 992 421439 1048
rect 413461 990 421439 992
rect 413461 987 413527 990
rect 421373 987 421439 990
rect 5257 914 5323 917
rect 11697 914 11763 917
rect 5257 912 11763 914
rect 5257 856 5262 912
rect 5318 856 11702 912
rect 11758 856 11763 912
rect 5257 854 11763 856
rect 5257 851 5323 854
rect 11697 851 11763 854
rect 19425 914 19491 917
rect 31017 914 31083 917
rect 19425 912 31083 914
rect 19425 856 19430 912
rect 19486 856 31022 912
rect 31078 856 31083 912
rect 19425 854 31083 856
rect 19425 851 19491 854
rect 31017 851 31083 854
rect 129365 914 129431 917
rect 140681 914 140747 917
rect 129365 912 140747 914
rect 129365 856 129370 912
rect 129426 856 140686 912
rect 140742 856 140747 912
rect 129365 854 140747 856
rect 129365 851 129431 854
rect 140681 851 140747 854
rect 181437 914 181503 917
rect 189257 914 189323 917
rect 181437 912 189323 914
rect 181437 856 181442 912
rect 181498 856 189262 912
rect 189318 856 189323 912
rect 181437 854 189323 856
rect 181437 851 181503 854
rect 189257 851 189323 854
rect 192017 914 192083 917
rect 199193 914 199259 917
rect 192017 912 199259 914
rect 192017 856 192022 912
rect 192078 856 199198 912
rect 199254 856 199259 912
rect 192017 854 199259 856
rect 192017 851 192083 854
rect 199193 851 199259 854
rect 331765 914 331831 917
rect 333881 914 333947 917
rect 331765 912 333947 914
rect 331765 856 331770 912
rect 331826 856 333886 912
rect 333942 856 333947 912
rect 331765 854 333947 856
rect 331765 851 331831 854
rect 333881 851 333947 854
rect 400121 914 400187 917
rect 412357 914 412423 917
rect 420177 914 420243 917
rect 400121 912 402990 914
rect 400121 856 400126 912
rect 400182 856 402990 912
rect 400121 854 402990 856
rect 400121 851 400187 854
rect 8753 778 8819 781
rect 17861 778 17927 781
rect 8753 776 17927 778
rect 8753 720 8758 776
rect 8814 720 17866 776
rect 17922 720 17927 776
rect 8753 718 17927 720
rect 8753 715 8819 718
rect 17861 715 17927 718
rect 18229 778 18295 781
rect 36905 778 36971 781
rect 102041 778 102107 781
rect 18229 776 36971 778
rect 18229 720 18234 776
rect 18290 720 36910 776
rect 36966 720 36971 776
rect 18229 718 36971 720
rect 18229 715 18295 718
rect 36905 715 36971 718
rect 97950 776 102107 778
rect 97950 720 102046 776
rect 102102 720 102107 776
rect 97950 718 102107 720
rect 4061 642 4127 645
rect 9581 642 9647 645
rect 4061 640 9647 642
rect 4061 584 4066 640
rect 4122 584 9586 640
rect 9642 584 9647 640
rect 4061 582 9647 584
rect 4061 579 4127 582
rect 9581 579 9647 582
rect 11145 642 11211 645
rect 28257 642 28323 645
rect 11145 640 28323 642
rect 11145 584 11150 640
rect 11206 584 28262 640
rect 28318 584 28323 640
rect 11145 582 28323 584
rect 11145 579 11211 582
rect 28257 579 28323 582
rect 31293 642 31359 645
rect 33225 642 33291 645
rect 31293 640 33291 642
rect 31293 584 31298 640
rect 31354 584 33230 640
rect 33286 584 33291 640
rect 31293 582 33291 584
rect 31293 579 31359 582
rect 33225 579 33291 582
rect 77385 642 77451 645
rect 92105 642 92171 645
rect 77385 640 92171 642
rect 77385 584 77390 640
rect 77446 584 92110 640
rect 92166 584 92171 640
rect 77385 582 92171 584
rect 77385 579 77451 582
rect 92105 579 92171 582
rect 8201 506 8267 509
rect 26969 506 27035 509
rect 8201 504 27035 506
rect 8201 448 8206 504
rect 8262 448 26974 504
rect 27030 448 27035 504
rect 8201 446 27035 448
rect 8201 443 8267 446
rect 26969 443 27035 446
rect 28165 506 28231 509
rect 36997 506 37063 509
rect 28165 504 37063 506
rect 28165 448 28170 504
rect 28226 448 37002 504
rect 37058 448 37063 504
rect 28165 446 37063 448
rect 28165 443 28231 446
rect 36997 443 37063 446
rect 83457 506 83523 509
rect 97625 506 97691 509
rect 83457 504 97691 506
rect 83457 448 83462 504
rect 83518 448 97630 504
rect 97686 448 97691 504
rect 83457 446 97691 448
rect 83457 443 83523 446
rect 97625 443 97691 446
rect 3325 370 3391 373
rect 22553 370 22619 373
rect 3325 368 22619 370
rect 3325 312 3330 368
rect 3386 312 22558 368
rect 22614 312 22619 368
rect 3325 310 22619 312
rect 3325 307 3391 310
rect 22553 307 22619 310
rect 24761 370 24827 373
rect 30281 370 30347 373
rect 24761 368 30347 370
rect 24761 312 24766 368
rect 24822 312 30286 368
rect 30342 312 30347 368
rect 24761 310 30347 312
rect 24761 307 24827 310
rect 30281 307 30347 310
rect 84653 370 84719 373
rect 87781 370 87847 373
rect 97950 370 98010 718
rect 102041 715 102107 718
rect 123477 778 123543 781
rect 135161 778 135227 781
rect 123477 776 135227 778
rect 123477 720 123482 776
rect 123538 720 135166 776
rect 135222 720 135227 776
rect 123477 718 135227 720
rect 123477 715 123543 718
rect 135161 715 135227 718
rect 136449 778 136515 781
rect 147305 778 147371 781
rect 136449 776 147371 778
rect 136449 720 136454 776
rect 136510 720 147310 776
rect 147366 720 147371 776
rect 136449 718 147371 720
rect 136449 715 136515 718
rect 147305 715 147371 718
rect 167177 778 167243 781
rect 176009 778 176075 781
rect 167177 776 176075 778
rect 167177 720 167182 776
rect 167238 720 176014 776
rect 176070 720 176075 776
rect 167177 718 176075 720
rect 167177 715 167243 718
rect 176009 715 176075 718
rect 179045 778 179111 781
rect 187049 778 187115 781
rect 179045 776 187115 778
rect 179045 720 179050 776
rect 179106 720 187054 776
rect 187110 720 187115 776
rect 179045 718 187115 720
rect 179045 715 179111 718
rect 187049 715 187115 718
rect 190821 778 190887 781
rect 198089 778 198155 781
rect 190821 776 198155 778
rect 190821 720 190826 776
rect 190882 720 198094 776
rect 198150 720 198155 776
rect 190821 718 198155 720
rect 190821 715 190887 718
rect 198089 715 198155 718
rect 199101 778 199167 781
rect 205817 778 205883 781
rect 199101 776 205883 778
rect 199101 720 199106 776
rect 199162 720 205822 776
rect 205878 720 205883 776
rect 199101 718 205883 720
rect 199101 715 199167 718
rect 205817 715 205883 718
rect 130561 642 130627 645
rect 132769 642 132835 645
rect 130561 640 132835 642
rect 130561 584 130566 640
rect 130622 584 132774 640
rect 132830 584 132835 640
rect 130561 582 132835 584
rect 130561 579 130627 582
rect 132769 579 132835 582
rect 132953 642 133019 645
rect 143993 642 144059 645
rect 132953 640 144059 642
rect 132953 584 132958 640
rect 133014 584 143998 640
rect 144054 584 144059 640
rect 132953 582 144059 584
rect 132953 579 133019 582
rect 143993 579 144059 582
rect 173157 642 173223 645
rect 181529 642 181595 645
rect 184841 642 184907 645
rect 195881 642 195947 645
rect 173157 640 181595 642
rect 173157 584 173162 640
rect 173218 584 181534 640
rect 181590 584 181595 640
rect 173157 582 181595 584
rect 173157 579 173223 582
rect 181529 579 181595 582
rect 182774 640 184907 642
rect 182774 584 184846 640
rect 184902 584 184907 640
rect 182774 582 184907 584
rect 98821 506 98887 509
rect 130745 506 130811 509
rect 98821 504 98930 506
rect 98821 448 98826 504
rect 98882 448 98930 504
rect 98821 443 98930 448
rect 84653 368 87706 370
rect 84653 312 84658 368
rect 84714 312 87706 368
rect 84653 310 87706 312
rect 84653 307 84719 310
rect 1485 234 1551 237
rect 21449 234 21515 237
rect 1485 232 21515 234
rect 1485 176 1490 232
rect 1546 176 21454 232
rect 21510 176 21515 232
rect 1485 174 21515 176
rect 1485 171 1551 174
rect 21449 171 21515 174
rect 26325 234 26391 237
rect 44633 234 44699 237
rect 26325 232 44699 234
rect 26325 176 26330 232
rect 26386 176 44638 232
rect 44694 176 44699 232
rect 26325 174 44699 176
rect 87646 234 87706 310
rect 87781 368 98010 370
rect 87781 312 87786 368
rect 87842 312 98010 368
rect 87781 310 98010 312
rect 87781 307 87847 310
rect 98870 234 98930 443
rect 87646 174 98930 234
rect 122790 504 130811 506
rect 122790 448 130750 504
rect 130806 448 130811 504
rect 122790 446 130811 448
rect 26325 171 26391 174
rect 44633 171 44699 174
rect 381 98 447 101
rect 20345 98 20411 101
rect 381 96 20411 98
rect 381 40 386 96
rect 442 40 20350 96
rect 20406 40 20411 96
rect 381 38 20411 40
rect 381 35 447 38
rect 20345 35 20411 38
rect 44633 98 44699 101
rect 61193 98 61259 101
rect 44633 96 61259 98
rect 44633 40 44638 96
rect 44694 40 61198 96
rect 61254 40 61259 96
rect 44633 38 61259 40
rect 44633 35 44699 38
rect 61193 35 61259 38
rect 90173 98 90239 101
rect 104157 98 104223 101
rect 90173 96 104223 98
rect 90173 40 90178 96
rect 90234 40 104162 96
rect 104218 40 104223 96
rect 90173 38 104223 40
rect 90173 35 90239 38
rect 104157 35 104223 38
rect 119153 98 119219 101
rect 122790 98 122850 446
rect 130745 443 130811 446
rect 148501 506 148567 509
rect 160277 506 160343 509
rect 169385 506 169451 509
rect 148501 504 148610 506
rect 148501 448 148506 504
rect 148562 448 148610 504
rect 148501 443 148610 448
rect 160277 504 169451 506
rect 160277 448 160282 504
rect 160338 448 169390 504
rect 169446 448 169451 504
rect 160277 446 169451 448
rect 160277 443 160343 446
rect 169385 443 169451 446
rect 170581 506 170647 509
rect 179321 506 179387 509
rect 170581 504 179387 506
rect 170581 448 170586 504
rect 170642 448 179326 504
rect 179382 448 179387 504
rect 170581 446 179387 448
rect 170581 443 170647 446
rect 179321 443 179387 446
rect 127157 370 127223 373
rect 138473 370 138539 373
rect 127157 368 138539 370
rect 127157 312 127162 368
rect 127218 312 138478 368
rect 138534 312 138539 368
rect 127157 310 138539 312
rect 127157 307 127223 310
rect 138473 307 138539 310
rect 125685 234 125751 237
rect 137277 234 137343 237
rect 125685 232 137343 234
rect 125685 176 125690 232
rect 125746 176 137282 232
rect 137338 176 137343 232
rect 125685 174 137343 176
rect 125685 171 125751 174
rect 137277 171 137343 174
rect 137461 234 137527 237
rect 148550 234 148610 443
rect 165889 370 165955 373
rect 174905 370 174971 373
rect 165889 368 174971 370
rect 165889 312 165894 368
rect 165950 312 174910 368
rect 174966 312 174971 368
rect 165889 310 174971 312
rect 165889 307 165955 310
rect 174905 307 174971 310
rect 176837 370 176903 373
rect 182774 370 182834 582
rect 184841 579 184907 582
rect 192710 640 195947 642
rect 192710 584 195886 640
rect 195942 584 195947 640
rect 192710 582 195947 584
rect 402930 642 402990 854
rect 412357 912 420243 914
rect 412357 856 412362 912
rect 412418 856 420182 912
rect 420238 856 420243 912
rect 412357 854 420243 856
rect 412357 851 412423 854
rect 420177 851 420243 854
rect 481909 914 481975 917
rect 494697 914 494763 917
rect 481909 912 494763 914
rect 481909 856 481914 912
rect 481970 856 494702 912
rect 494758 856 494763 912
rect 481909 854 494763 856
rect 481909 851 481975 854
rect 494697 851 494763 854
rect 552565 914 552631 917
rect 570321 914 570387 917
rect 552565 912 570387 914
rect 552565 856 552570 912
rect 552626 856 570326 912
rect 570382 856 570387 912
rect 552565 854 570387 856
rect 552565 851 552631 854
rect 570321 851 570387 854
rect 417877 778 417943 781
rect 426157 778 426223 781
rect 417877 776 426223 778
rect 417877 720 417882 776
rect 417938 720 426162 776
rect 426218 720 426223 776
rect 417877 718 426223 720
rect 417877 715 417943 718
rect 426157 715 426223 718
rect 475285 778 475351 781
rect 487613 778 487679 781
rect 475285 776 487679 778
rect 475285 720 475290 776
rect 475346 720 487618 776
rect 487674 720 487679 776
rect 475285 718 487679 720
rect 475285 715 475351 718
rect 487613 715 487679 718
rect 534901 778 534967 781
rect 545941 778 546007 781
rect 563237 778 563303 781
rect 534901 776 538230 778
rect 534901 720 534906 776
rect 534962 720 538230 776
rect 534901 718 538230 720
rect 534901 715 534967 718
rect 407205 642 407271 645
rect 402930 640 407271 642
rect 402930 584 407210 640
rect 407266 584 407271 640
rect 402930 582 407271 584
rect 176837 368 182834 370
rect 176837 312 176842 368
rect 176898 312 182834 368
rect 176837 310 182834 312
rect 188981 370 189047 373
rect 192710 370 192770 582
rect 195881 579 195947 582
rect 407205 579 407271 582
rect 411161 642 411227 645
rect 418981 642 419047 645
rect 411161 640 419047 642
rect 411161 584 411166 640
rect 411222 584 418986 640
rect 419042 584 419047 640
rect 411161 582 419047 584
rect 411161 579 411227 582
rect 418981 579 419047 582
rect 420085 642 420151 645
rect 428457 642 428523 645
rect 420085 640 428523 642
rect 420085 584 420090 640
rect 420146 584 428462 640
rect 428518 584 428523 640
rect 420085 582 428523 584
rect 420085 579 420151 582
rect 428457 579 428523 582
rect 480805 642 480871 645
rect 493501 642 493567 645
rect 480805 640 493567 642
rect 480805 584 480810 640
rect 480866 584 493506 640
rect 493562 584 493567 640
rect 480805 582 493567 584
rect 480805 579 480871 582
rect 493501 579 493567 582
rect 498469 642 498535 645
rect 512453 642 512519 645
rect 517145 642 517211 645
rect 498469 640 512519 642
rect 498469 584 498474 640
rect 498530 584 512458 640
rect 512514 584 512519 640
rect 498469 582 512519 584
rect 498469 579 498535 582
rect 512453 579 512519 582
rect 515630 640 517211 642
rect 515630 584 517150 640
rect 517206 584 517211 640
rect 515630 582 517211 584
rect 414565 506 414631 509
rect 447685 506 447751 509
rect 457713 506 457779 509
rect 414565 504 422310 506
rect 414565 448 414570 504
rect 414626 448 422310 504
rect 414565 446 422310 448
rect 414565 443 414631 446
rect 188981 368 192770 370
rect 188981 312 188986 368
rect 189042 312 192770 368
rect 188981 310 192770 312
rect 198365 370 198431 373
rect 204713 370 204779 373
rect 198365 368 204779 370
rect 198365 312 198370 368
rect 198426 312 204718 368
rect 204774 312 204779 368
rect 198365 310 204779 312
rect 176837 307 176903 310
rect 188981 307 189047 310
rect 198365 307 198431 310
rect 204713 307 204779 310
rect 405641 370 405707 373
rect 412817 370 412883 373
rect 405641 368 412883 370
rect 405641 312 405646 368
rect 405702 312 412822 368
rect 412878 312 412883 368
rect 405641 310 412883 312
rect 422250 370 422310 446
rect 447685 504 457779 506
rect 447685 448 447690 504
rect 447746 448 457718 504
rect 457774 448 457779 504
rect 447685 446 457779 448
rect 447685 443 447751 446
rect 457713 443 457779 446
rect 465349 506 465415 509
rect 476389 506 476455 509
rect 465349 504 476455 506
rect 465349 448 465354 504
rect 465410 448 476394 504
rect 476450 448 476455 504
rect 465349 446 476455 448
rect 465349 443 465415 446
rect 476389 443 476455 446
rect 478597 506 478663 509
rect 490741 506 490807 509
rect 478597 504 490807 506
rect 478597 448 478602 504
rect 478658 448 490746 504
rect 490802 448 490807 504
rect 478597 446 490807 448
rect 478597 443 478663 446
rect 490741 443 490807 446
rect 492949 506 493015 509
rect 506657 506 506723 509
rect 492949 504 506723 506
rect 492949 448 492954 504
rect 493010 448 506662 504
rect 506718 448 506723 504
rect 492949 446 506723 448
rect 492949 443 493015 446
rect 506657 443 506723 446
rect 422753 370 422819 373
rect 422250 368 422819 370
rect 422250 312 422758 368
rect 422814 312 422819 368
rect 422250 310 422819 312
rect 405641 307 405707 310
rect 412817 307 412883 310
rect 422753 307 422819 310
rect 428917 370 428983 373
rect 437473 370 437539 373
rect 428917 368 437539 370
rect 428917 312 428922 368
rect 428978 312 437478 368
rect 437534 312 437539 368
rect 428917 310 437539 312
rect 428917 307 428983 310
rect 437473 307 437539 310
rect 486141 370 486207 373
rect 498929 370 498995 373
rect 486141 368 498995 370
rect 486141 312 486146 368
rect 486202 312 498934 368
rect 498990 312 498995 368
rect 486141 310 498995 312
rect 486141 307 486207 310
rect 498929 307 498995 310
rect 502057 370 502123 373
rect 515489 370 515555 373
rect 502057 368 515555 370
rect 502057 312 502062 368
rect 502118 312 515494 368
rect 515550 312 515555 368
rect 502057 310 515555 312
rect 502057 307 502123 310
rect 515489 307 515555 310
rect 137461 232 148610 234
rect 137461 176 137466 232
rect 137522 176 148610 232
rect 137461 174 148610 176
rect 182357 234 182423 237
rect 190361 234 190427 237
rect 182357 232 190427 234
rect 182357 176 182362 232
rect 182418 176 190366 232
rect 190422 176 190427 232
rect 182357 174 190427 176
rect 137461 171 137527 174
rect 182357 171 182423 174
rect 190361 171 190427 174
rect 426709 234 426775 237
rect 435357 234 435423 237
rect 426709 232 435423 234
rect 426709 176 426714 232
rect 426770 176 435362 232
rect 435418 176 435423 232
rect 426709 174 435423 176
rect 426709 171 426775 174
rect 435357 171 435423 174
rect 487245 234 487311 237
rect 500309 234 500375 237
rect 487245 232 500375 234
rect 487245 176 487250 232
rect 487306 176 500314 232
rect 500370 176 500375 232
rect 487245 174 500375 176
rect 487245 171 487311 174
rect 500309 171 500375 174
rect 502701 234 502767 237
rect 515630 234 515690 582
rect 517145 579 517211 582
rect 519353 506 519419 509
rect 502701 232 515690 234
rect 502701 176 502706 232
rect 502762 176 515690 232
rect 502701 174 515690 176
rect 519310 504 519419 506
rect 519310 448 519358 504
rect 519414 448 519419 504
rect 519310 443 519419 448
rect 502701 171 502767 174
rect 119153 96 122850 98
rect 119153 40 119158 96
rect 119214 40 122850 96
rect 119153 38 122850 40
rect 139853 98 139919 101
rect 150341 98 150407 101
rect 139853 96 150407 98
rect 139853 40 139858 96
rect 139914 40 150346 96
rect 150402 40 150407 96
rect 139853 38 150407 40
rect 119153 35 119219 38
rect 139853 35 139919 38
rect 150341 35 150407 38
rect 159265 98 159331 101
rect 168005 98 168071 101
rect 159265 96 168071 98
rect 159265 40 159270 96
rect 159326 40 168010 96
rect 168066 40 168071 96
rect 159265 38 168071 40
rect 159265 35 159331 38
rect 168005 35 168071 38
rect 175825 98 175891 101
rect 183461 98 183527 101
rect 175825 96 183527 98
rect 175825 40 175830 96
rect 175886 40 183466 96
rect 183522 40 183527 96
rect 175825 38 183527 40
rect 175825 35 175891 38
rect 183461 35 183527 38
rect 187141 98 187207 101
rect 194777 98 194843 101
rect 187141 96 194843 98
rect 187141 40 187146 96
rect 187202 40 194782 96
rect 194838 40 194843 96
rect 187141 38 194843 40
rect 187141 35 187207 38
rect 194777 35 194843 38
rect 197169 98 197235 101
rect 203517 98 203583 101
rect 197169 96 203583 98
rect 197169 40 197174 96
rect 197230 40 203522 96
rect 203578 40 203583 96
rect 197169 38 203583 40
rect 197169 35 197235 38
rect 203517 35 203583 38
rect 390277 98 390343 101
rect 396165 98 396231 101
rect 390277 96 396231 98
rect 390277 40 390282 96
rect 390338 40 396170 96
rect 396226 40 396231 96
rect 390277 38 396231 40
rect 390277 35 390343 38
rect 396165 35 396231 38
rect 407941 98 408007 101
rect 415301 98 415367 101
rect 407941 96 415367 98
rect 407941 40 407946 96
rect 408002 40 415306 96
rect 415362 40 415367 96
rect 407941 38 415367 40
rect 407941 35 408007 38
rect 415301 35 415367 38
rect 457621 98 457687 101
rect 468477 98 468543 101
rect 457621 96 468543 98
rect 457621 40 457626 96
rect 457682 40 468482 96
rect 468538 40 468543 96
rect 457621 38 468543 40
rect 457621 35 457687 38
rect 468477 35 468543 38
rect 476297 98 476363 101
rect 488993 98 489059 101
rect 476297 96 489059 98
rect 476297 40 476302 96
rect 476358 40 488998 96
rect 489054 40 489059 96
rect 476297 38 489059 40
rect 476297 35 476363 38
rect 488993 35 489059 38
rect 489637 98 489703 101
rect 503161 98 503227 101
rect 489637 96 503227 98
rect 489637 40 489642 96
rect 489698 40 503166 96
rect 503222 40 503227 96
rect 489637 38 503227 40
rect 489637 35 489703 38
rect 503161 35 503227 38
rect 503713 98 503779 101
rect 518157 98 518223 101
rect 503713 96 518223 98
rect 503713 40 503718 96
rect 503774 40 518162 96
rect 518218 40 518223 96
rect 503713 38 518223 40
rect 519310 98 519370 443
rect 538170 370 538230 718
rect 545941 776 563303 778
rect 545941 720 545946 776
rect 546002 720 563242 776
rect 563298 720 563303 776
rect 545941 718 563303 720
rect 545941 715 546007 718
rect 563237 715 563303 718
rect 551369 642 551435 645
rect 569125 642 569191 645
rect 551369 640 569191 642
rect 551369 584 551374 640
rect 551430 584 569130 640
rect 569186 584 569191 640
rect 551369 582 569191 584
rect 551369 579 551435 582
rect 569125 579 569191 582
rect 559189 506 559255 509
rect 577129 506 577195 509
rect 559189 504 577195 506
rect 559189 448 559194 504
rect 559250 448 577134 504
rect 577190 448 577195 504
rect 559189 446 577195 448
rect 559189 443 559255 446
rect 577129 443 577195 446
rect 551645 370 551711 373
rect 538170 368 551711 370
rect 538170 312 551650 368
rect 551706 312 551711 368
rect 538170 310 551711 312
rect 551645 307 551711 310
rect 558085 370 558151 373
rect 575749 370 575815 373
rect 558085 368 575815 370
rect 558085 312 558090 368
rect 558146 312 575754 368
rect 575810 312 575815 368
rect 558085 310 575815 312
rect 558085 307 558151 310
rect 575749 307 575815 310
rect 526069 234 526135 237
rect 542169 234 542235 237
rect 526069 232 542235 234
rect 526069 176 526074 232
rect 526130 176 542174 232
rect 542230 176 542235 232
rect 526069 174 542235 176
rect 526069 171 526135 174
rect 542169 171 542235 174
rect 562501 234 562567 237
rect 581821 234 581887 237
rect 562501 232 581887 234
rect 562501 176 562506 232
rect 562562 176 581826 232
rect 581882 176 581887 232
rect 562501 174 581887 176
rect 562501 171 562567 174
rect 581821 171 581887 174
rect 534717 98 534783 101
rect 519310 96 534783 98
rect 519310 40 534722 96
rect 534778 40 534783 96
rect 519310 38 534783 40
rect 503713 35 503779 38
rect 518157 35 518223 38
rect 534717 35 534783 38
rect 544837 98 544903 101
rect 562225 98 562291 101
rect 544837 96 562291 98
rect 544837 40 544842 96
rect 544898 40 562230 96
rect 562286 40 562291 96
rect 544837 38 562291 40
rect 544837 35 544903 38
rect 562225 35 562291 38
rect 563605 98 563671 101
rect 583569 98 583635 101
rect 563605 96 583635 98
rect 563605 40 563610 96
rect 563666 40 583574 96
rect 583630 40 583635 96
rect 563605 38 583635 40
rect 563605 35 563671 38
rect 583569 35 583635 38
<< via3 >>
rect 3740 371316 3804 371380
rect 3556 358396 3620 358460
rect 3372 345340 3436 345404
rect 3740 344660 3804 344724
rect 574692 344660 574756 344724
rect 3556 330244 3620 330308
rect 574876 330244 574940 330308
rect 574692 325212 574756 325276
rect 3740 319228 3804 319292
rect 3372 315828 3436 315892
rect 575060 315828 575124 315892
rect 574876 312020 574940 312084
rect 3556 306172 3620 306236
rect 3740 301412 3804 301476
rect 574692 301412 574756 301476
rect 575060 298692 575124 298756
rect 3372 293116 3436 293180
rect 3556 286996 3620 287060
rect 575060 286996 575124 287060
rect 3372 272580 3436 272644
rect 574876 272580 574940 272644
rect 574692 272172 574756 272236
rect 8156 267140 8220 267204
rect 575060 258844 575124 258908
rect 8156 258164 8220 258228
rect 574692 258164 574756 258228
rect 7420 254084 7484 254148
rect 574876 245516 574940 245580
rect 7420 243748 7484 243812
rect 574876 243748 574940 243812
rect 7420 241028 7484 241092
rect 574692 232324 574756 232388
rect 7420 229332 7484 229396
rect 574692 229332 574756 229396
rect 574876 218996 574940 219060
rect 574876 214916 574940 214980
rect 574692 205668 574756 205732
rect 574692 200500 574756 200564
rect 574876 192476 574940 192540
rect 6316 188804 6380 188868
rect 6316 186084 6380 186148
rect 574876 186084 574940 186148
rect 574692 179148 574756 179212
rect 6316 171668 6380 171732
rect 574692 171668 574756 171732
rect 574876 165820 574940 165884
rect 6316 162828 6380 162892
rect 6316 157252 6380 157316
rect 574876 157252 574940 157316
rect 574692 152628 574756 152692
rect 6316 149772 6380 149836
rect 4844 142836 4908 142900
rect 574692 142836 574756 142900
rect 574876 139300 574940 139364
rect 4844 136716 4908 136780
rect 3372 128420 3436 128484
rect 574876 128420 574940 128484
rect 574692 125972 574756 126036
rect 3556 114004 3620 114068
rect 574692 114004 574756 114068
rect 574876 112780 574940 112844
rect 3372 110604 3436 110668
rect 8892 99588 8956 99652
rect 574876 99588 574940 99652
rect 574692 99452 574756 99516
rect 3556 97548 3620 97612
rect 574876 86124 574940 86188
rect 8708 85172 8772 85236
rect 574692 85172 574756 85236
rect 8892 84628 8956 84692
rect 574692 72932 574756 72996
rect 8708 71572 8772 71636
rect 8892 70756 8956 70820
rect 574692 70756 574756 70820
rect 574692 59604 574756 59668
rect 8892 58516 8956 58580
rect 8892 56340 8956 56404
rect 574692 56340 574756 56404
rect 574692 46276 574756 46340
rect 8892 45460 8956 45524
rect 8892 41924 8956 41988
rect 574692 41924 574756 41988
rect 574692 33084 574756 33148
rect 8892 32404 8956 32468
rect 6316 27508 6380 27572
rect 575428 27508 575492 27572
rect 575428 19756 575492 19820
rect 6316 19348 6380 19412
rect 8892 13092 8956 13156
rect 574692 13092 574756 13156
rect 574692 6564 574756 6628
rect 8892 6428 8956 6492
rect 47900 3844 47964 3908
rect 59860 3844 59924 3908
rect 383516 3708 383580 3772
rect 389404 3708 389468 3772
rect 533476 3708 533540 3772
rect 34836 3164 34900 3228
rect 47900 2680 47964 2684
rect 47900 2624 47914 2680
rect 47914 2624 47964 2680
rect 47900 2620 47964 2624
rect 34836 2544 34900 2548
rect 34836 2488 34850 2544
rect 34850 2488 34900 2544
rect 34836 2484 34900 2488
rect 59860 2756 59924 2820
rect 364196 3028 364260 3092
rect 364196 2756 364260 2820
rect 377444 3028 377508 3092
rect 397500 3300 397564 3364
rect 405964 3164 406028 3228
rect 397500 2680 397564 2684
rect 397500 2624 397550 2680
rect 397550 2624 397564 2680
rect 397500 2620 397564 2624
rect 377444 2544 377508 2548
rect 377444 2488 377494 2544
rect 377494 2488 377508 2544
rect 377444 2484 377508 2488
rect 383516 2544 383580 2548
rect 383516 2488 383566 2544
rect 383566 2488 383580 2544
rect 383516 2484 383580 2488
rect 389404 2544 389468 2548
rect 405964 2816 406028 2820
rect 405964 2760 406014 2816
rect 406014 2760 406028 2816
rect 405964 2756 406028 2760
rect 462636 3572 462700 3636
rect 389404 2488 389454 2544
rect 389454 2488 389468 2544
rect 389404 2484 389468 2488
rect 463740 3436 463804 3500
rect 458404 3300 458468 3364
rect 467236 3300 467300 3364
rect 466316 3164 466380 3228
rect 458404 2892 458468 2956
rect 462636 2680 462700 2684
rect 463740 2756 463804 2820
rect 498148 3028 498212 3092
rect 462636 2624 462686 2680
rect 462686 2624 462700 2680
rect 462636 2620 462700 2624
rect 517836 3572 517900 3636
rect 526300 3572 526364 3636
rect 516732 3436 516796 3500
rect 514524 3164 514588 3228
rect 514524 2756 514588 2820
rect 516732 2892 516796 2956
rect 517836 3028 517900 3092
rect 522988 3028 523052 3092
rect 529980 3164 530044 3228
rect 526484 3028 526548 3092
rect 527588 3028 527652 3092
rect 526300 2892 526364 2956
rect 545252 3572 545316 3636
rect 533476 2892 533540 2956
rect 547644 3436 547708 3500
rect 552428 3300 552492 3364
rect 558500 3844 558564 3908
rect 533292 2756 533356 2820
rect 526484 2680 526548 2684
rect 526484 2624 526534 2680
rect 526534 2624 526548 2680
rect 526484 2620 526548 2624
rect 527588 2680 527652 2684
rect 527588 2624 527638 2680
rect 527638 2624 527652 2680
rect 527588 2620 527652 2624
rect 529980 2680 530044 2684
rect 529980 2624 530030 2680
rect 530030 2624 530044 2680
rect 529980 2620 530044 2624
rect 533292 2680 533356 2684
rect 533292 2624 533342 2680
rect 533342 2624 533356 2680
rect 533292 2620 533356 2624
rect 552428 2680 552492 2684
rect 552428 2624 552478 2680
rect 552478 2624 552492 2680
rect 552428 2620 552492 2624
rect 466316 2544 466380 2548
rect 466316 2488 466330 2544
rect 466330 2488 466380 2544
rect 466316 2484 466380 2488
rect 467236 2544 467300 2548
rect 467236 2488 467286 2544
rect 467286 2488 467300 2544
rect 467236 2484 467300 2488
rect 498148 2544 498212 2548
rect 498148 2488 498198 2544
rect 498198 2488 498212 2544
rect 498148 2484 498212 2488
rect 522988 2544 523052 2548
rect 522988 2488 523038 2544
rect 523038 2488 523052 2544
rect 522988 2484 523052 2488
rect 545252 2544 545316 2548
rect 545252 2488 545302 2544
rect 545302 2488 545316 2544
rect 545252 2484 545316 2488
rect 547644 2484 547708 2548
rect 558500 2816 558564 2820
rect 558500 2760 558550 2816
rect 558550 2760 558564 2816
rect 558500 2756 558564 2760
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711002 -8694 711558
rect -8138 711002 -8106 711558
rect -8726 677494 -8106 711002
rect -8726 676938 -8694 677494
rect -8138 676938 -8106 677494
rect -8726 641494 -8106 676938
rect -8726 640938 -8694 641494
rect -8138 640938 -8106 641494
rect -8726 605494 -8106 640938
rect -8726 604938 -8694 605494
rect -8138 604938 -8106 605494
rect -8726 569494 -8106 604938
rect -8726 568938 -8694 569494
rect -8138 568938 -8106 569494
rect -8726 533494 -8106 568938
rect -8726 532938 -8694 533494
rect -8138 532938 -8106 533494
rect -8726 497494 -8106 532938
rect -8726 496938 -8694 497494
rect -8138 496938 -8106 497494
rect -8726 461494 -8106 496938
rect -8726 460938 -8694 461494
rect -8138 460938 -8106 461494
rect -8726 425494 -8106 460938
rect -8726 424938 -8694 425494
rect -8138 424938 -8106 425494
rect -8726 389494 -8106 424938
rect -8726 388938 -8694 389494
rect -8138 388938 -8106 389494
rect -8726 353494 -8106 388938
rect -8726 352938 -8694 353494
rect -8138 352938 -8106 353494
rect -8726 317494 -8106 352938
rect -8726 316938 -8694 317494
rect -8138 316938 -8106 317494
rect -8726 281494 -8106 316938
rect -8726 280938 -8694 281494
rect -8138 280938 -8106 281494
rect -8726 245494 -8106 280938
rect -8726 244938 -8694 245494
rect -8138 244938 -8106 245494
rect -8726 209494 -8106 244938
rect -8726 208938 -8694 209494
rect -8138 208938 -8106 209494
rect -8726 173494 -8106 208938
rect -8726 172938 -8694 173494
rect -8138 172938 -8106 173494
rect -8726 137494 -8106 172938
rect -8726 136938 -8694 137494
rect -8138 136938 -8106 137494
rect -8726 101494 -8106 136938
rect -8726 100938 -8694 101494
rect -8138 100938 -8106 101494
rect -8726 65494 -8106 100938
rect -8726 64938 -8694 65494
rect -8138 64938 -8106 65494
rect -8726 29494 -8106 64938
rect -8726 28938 -8694 29494
rect -8138 28938 -8106 29494
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710042 -7734 710598
rect -7178 710042 -7146 710598
rect -7766 673774 -7146 710042
rect -7766 673218 -7734 673774
rect -7178 673218 -7146 673774
rect -7766 637774 -7146 673218
rect -7766 637218 -7734 637774
rect -7178 637218 -7146 637774
rect -7766 601774 -7146 637218
rect -7766 601218 -7734 601774
rect -7178 601218 -7146 601774
rect -7766 565774 -7146 601218
rect -7766 565218 -7734 565774
rect -7178 565218 -7146 565774
rect -7766 529774 -7146 565218
rect -7766 529218 -7734 529774
rect -7178 529218 -7146 529774
rect -7766 493774 -7146 529218
rect -7766 493218 -7734 493774
rect -7178 493218 -7146 493774
rect -7766 457774 -7146 493218
rect -7766 457218 -7734 457774
rect -7178 457218 -7146 457774
rect -7766 421774 -7146 457218
rect -7766 421218 -7734 421774
rect -7178 421218 -7146 421774
rect -7766 385774 -7146 421218
rect -7766 385218 -7734 385774
rect -7178 385218 -7146 385774
rect -7766 349774 -7146 385218
rect -7766 349218 -7734 349774
rect -7178 349218 -7146 349774
rect -7766 313774 -7146 349218
rect -7766 313218 -7734 313774
rect -7178 313218 -7146 313774
rect -7766 277774 -7146 313218
rect -7766 277218 -7734 277774
rect -7178 277218 -7146 277774
rect -7766 241774 -7146 277218
rect -7766 241218 -7734 241774
rect -7178 241218 -7146 241774
rect -7766 205774 -7146 241218
rect -7766 205218 -7734 205774
rect -7178 205218 -7146 205774
rect -7766 169774 -7146 205218
rect -7766 169218 -7734 169774
rect -7178 169218 -7146 169774
rect -7766 133774 -7146 169218
rect -7766 133218 -7734 133774
rect -7178 133218 -7146 133774
rect -7766 97774 -7146 133218
rect -7766 97218 -7734 97774
rect -7178 97218 -7146 97774
rect -7766 61774 -7146 97218
rect -7766 61218 -7734 61774
rect -7178 61218 -7146 61774
rect -7766 25774 -7146 61218
rect -7766 25218 -7734 25774
rect -7178 25218 -7146 25774
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709082 -6774 709638
rect -6218 709082 -6186 709638
rect -6806 670054 -6186 709082
rect -6806 669498 -6774 670054
rect -6218 669498 -6186 670054
rect -6806 634054 -6186 669498
rect -6806 633498 -6774 634054
rect -6218 633498 -6186 634054
rect -6806 598054 -6186 633498
rect -6806 597498 -6774 598054
rect -6218 597498 -6186 598054
rect -6806 562054 -6186 597498
rect -6806 561498 -6774 562054
rect -6218 561498 -6186 562054
rect -6806 526054 -6186 561498
rect -6806 525498 -6774 526054
rect -6218 525498 -6186 526054
rect -6806 490054 -6186 525498
rect -6806 489498 -6774 490054
rect -6218 489498 -6186 490054
rect -6806 454054 -6186 489498
rect -6806 453498 -6774 454054
rect -6218 453498 -6186 454054
rect -6806 418054 -6186 453498
rect -6806 417498 -6774 418054
rect -6218 417498 -6186 418054
rect -6806 382054 -6186 417498
rect -6806 381498 -6774 382054
rect -6218 381498 -6186 382054
rect -6806 346054 -6186 381498
rect -6806 345498 -6774 346054
rect -6218 345498 -6186 346054
rect -6806 310054 -6186 345498
rect -6806 309498 -6774 310054
rect -6218 309498 -6186 310054
rect -6806 274054 -6186 309498
rect -6806 273498 -6774 274054
rect -6218 273498 -6186 274054
rect -6806 238054 -6186 273498
rect -6806 237498 -6774 238054
rect -6218 237498 -6186 238054
rect -6806 202054 -6186 237498
rect -6806 201498 -6774 202054
rect -6218 201498 -6186 202054
rect -6806 166054 -6186 201498
rect -6806 165498 -6774 166054
rect -6218 165498 -6186 166054
rect -6806 130054 -6186 165498
rect -6806 129498 -6774 130054
rect -6218 129498 -6186 130054
rect -6806 94054 -6186 129498
rect -6806 93498 -6774 94054
rect -6218 93498 -6186 94054
rect -6806 58054 -6186 93498
rect -6806 57498 -6774 58054
rect -6218 57498 -6186 58054
rect -6806 22054 -6186 57498
rect -6806 21498 -6774 22054
rect -6218 21498 -6186 22054
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708122 -5814 708678
rect -5258 708122 -5226 708678
rect -5846 666334 -5226 708122
rect -5846 665778 -5814 666334
rect -5258 665778 -5226 666334
rect -5846 630334 -5226 665778
rect -5846 629778 -5814 630334
rect -5258 629778 -5226 630334
rect -5846 594334 -5226 629778
rect -5846 593778 -5814 594334
rect -5258 593778 -5226 594334
rect -5846 558334 -5226 593778
rect -5846 557778 -5814 558334
rect -5258 557778 -5226 558334
rect -5846 522334 -5226 557778
rect -5846 521778 -5814 522334
rect -5258 521778 -5226 522334
rect -5846 486334 -5226 521778
rect -5846 485778 -5814 486334
rect -5258 485778 -5226 486334
rect -5846 450334 -5226 485778
rect -5846 449778 -5814 450334
rect -5258 449778 -5226 450334
rect -5846 414334 -5226 449778
rect -5846 413778 -5814 414334
rect -5258 413778 -5226 414334
rect -5846 378334 -5226 413778
rect -5846 377778 -5814 378334
rect -5258 377778 -5226 378334
rect -5846 342334 -5226 377778
rect -5846 341778 -5814 342334
rect -5258 341778 -5226 342334
rect -5846 306334 -5226 341778
rect -5846 305778 -5814 306334
rect -5258 305778 -5226 306334
rect -5846 270334 -5226 305778
rect -5846 269778 -5814 270334
rect -5258 269778 -5226 270334
rect -5846 234334 -5226 269778
rect -5846 233778 -5814 234334
rect -5258 233778 -5226 234334
rect -5846 198334 -5226 233778
rect -5846 197778 -5814 198334
rect -5258 197778 -5226 198334
rect -5846 162334 -5226 197778
rect -5846 161778 -5814 162334
rect -5258 161778 -5226 162334
rect -5846 126334 -5226 161778
rect -5846 125778 -5814 126334
rect -5258 125778 -5226 126334
rect -5846 90334 -5226 125778
rect -5846 89778 -5814 90334
rect -5258 89778 -5226 90334
rect -5846 54334 -5226 89778
rect -5846 53778 -5814 54334
rect -5258 53778 -5226 54334
rect -5846 18334 -5226 53778
rect -5846 17778 -5814 18334
rect -5258 17778 -5226 18334
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707162 -4854 707718
rect -4298 707162 -4266 707718
rect -4886 698614 -4266 707162
rect -4886 698058 -4854 698614
rect -4298 698058 -4266 698614
rect -4886 662614 -4266 698058
rect -4886 662058 -4854 662614
rect -4298 662058 -4266 662614
rect -4886 626614 -4266 662058
rect -4886 626058 -4854 626614
rect -4298 626058 -4266 626614
rect -4886 590614 -4266 626058
rect -4886 590058 -4854 590614
rect -4298 590058 -4266 590614
rect -4886 554614 -4266 590058
rect -4886 554058 -4854 554614
rect -4298 554058 -4266 554614
rect -4886 518614 -4266 554058
rect -4886 518058 -4854 518614
rect -4298 518058 -4266 518614
rect -4886 482614 -4266 518058
rect -4886 482058 -4854 482614
rect -4298 482058 -4266 482614
rect -4886 446614 -4266 482058
rect -4886 446058 -4854 446614
rect -4298 446058 -4266 446614
rect -4886 410614 -4266 446058
rect -4886 410058 -4854 410614
rect -4298 410058 -4266 410614
rect -4886 374614 -4266 410058
rect -4886 374058 -4854 374614
rect -4298 374058 -4266 374614
rect -4886 338614 -4266 374058
rect -4886 338058 -4854 338614
rect -4298 338058 -4266 338614
rect -4886 302614 -4266 338058
rect -4886 302058 -4854 302614
rect -4298 302058 -4266 302614
rect -4886 266614 -4266 302058
rect -4886 266058 -4854 266614
rect -4298 266058 -4266 266614
rect -4886 230614 -4266 266058
rect -4886 230058 -4854 230614
rect -4298 230058 -4266 230614
rect -4886 194614 -4266 230058
rect -4886 194058 -4854 194614
rect -4298 194058 -4266 194614
rect -4886 158614 -4266 194058
rect -4886 158058 -4854 158614
rect -4298 158058 -4266 158614
rect -4886 122614 -4266 158058
rect -4886 122058 -4854 122614
rect -4298 122058 -4266 122614
rect -4886 86614 -4266 122058
rect -4886 86058 -4854 86614
rect -4298 86058 -4266 86614
rect -4886 50614 -4266 86058
rect -4886 50058 -4854 50614
rect -4298 50058 -4266 50614
rect -4886 14614 -4266 50058
rect -4886 14058 -4854 14614
rect -4298 14058 -4266 14614
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706202 -3894 706758
rect -3338 706202 -3306 706758
rect -3926 694894 -3306 706202
rect -3926 694338 -3894 694894
rect -3338 694338 -3306 694894
rect -3926 658894 -3306 694338
rect -3926 658338 -3894 658894
rect -3338 658338 -3306 658894
rect -3926 622894 -3306 658338
rect -3926 622338 -3894 622894
rect -3338 622338 -3306 622894
rect -3926 586894 -3306 622338
rect -3926 586338 -3894 586894
rect -3338 586338 -3306 586894
rect -3926 550894 -3306 586338
rect -3926 550338 -3894 550894
rect -3338 550338 -3306 550894
rect -3926 514894 -3306 550338
rect -3926 514338 -3894 514894
rect -3338 514338 -3306 514894
rect -3926 478894 -3306 514338
rect -3926 478338 -3894 478894
rect -3338 478338 -3306 478894
rect -3926 442894 -3306 478338
rect -3926 442338 -3894 442894
rect -3338 442338 -3306 442894
rect -3926 406894 -3306 442338
rect -3926 406338 -3894 406894
rect -3338 406338 -3306 406894
rect -3926 370894 -3306 406338
rect -3926 370338 -3894 370894
rect -3338 370338 -3306 370894
rect -3926 334894 -3306 370338
rect -3926 334338 -3894 334894
rect -3338 334338 -3306 334894
rect -3926 298894 -3306 334338
rect -3926 298338 -3894 298894
rect -3338 298338 -3306 298894
rect -3926 262894 -3306 298338
rect -3926 262338 -3894 262894
rect -3338 262338 -3306 262894
rect -3926 226894 -3306 262338
rect -3926 226338 -3894 226894
rect -3338 226338 -3306 226894
rect -3926 190894 -3306 226338
rect -3926 190338 -3894 190894
rect -3338 190338 -3306 190894
rect -3926 154894 -3306 190338
rect -3926 154338 -3894 154894
rect -3338 154338 -3306 154894
rect -3926 118894 -3306 154338
rect -3926 118338 -3894 118894
rect -3338 118338 -3306 118894
rect -3926 82894 -3306 118338
rect -3926 82338 -3894 82894
rect -3338 82338 -3306 82894
rect -3926 46894 -3306 82338
rect -3926 46338 -3894 46894
rect -3338 46338 -3306 46894
rect -3926 10894 -3306 46338
rect -3926 10338 -3894 10894
rect -3338 10338 -3306 10894
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705242 -2934 705798
rect -2378 705242 -2346 705798
rect -2966 691174 -2346 705242
rect -2966 690618 -2934 691174
rect -2378 690618 -2346 691174
rect -2966 655174 -2346 690618
rect -2966 654618 -2934 655174
rect -2378 654618 -2346 655174
rect -2966 619174 -2346 654618
rect -2966 618618 -2934 619174
rect -2378 618618 -2346 619174
rect -2966 583174 -2346 618618
rect -2966 582618 -2934 583174
rect -2378 582618 -2346 583174
rect -2966 547174 -2346 582618
rect -2966 546618 -2934 547174
rect -2378 546618 -2346 547174
rect -2966 511174 -2346 546618
rect -2966 510618 -2934 511174
rect -2378 510618 -2346 511174
rect -2966 475174 -2346 510618
rect -2966 474618 -2934 475174
rect -2378 474618 -2346 475174
rect -2966 439174 -2346 474618
rect -2966 438618 -2934 439174
rect -2378 438618 -2346 439174
rect -2966 403174 -2346 438618
rect -2966 402618 -2934 403174
rect -2378 402618 -2346 403174
rect -2966 367174 -2346 402618
rect -2966 366618 -2934 367174
rect -2378 366618 -2346 367174
rect -2966 331174 -2346 366618
rect -2966 330618 -2934 331174
rect -2378 330618 -2346 331174
rect -2966 295174 -2346 330618
rect -2966 294618 -2934 295174
rect -2378 294618 -2346 295174
rect -2966 259174 -2346 294618
rect -2966 258618 -2934 259174
rect -2378 258618 -2346 259174
rect -2966 223174 -2346 258618
rect -2966 222618 -2934 223174
rect -2378 222618 -2346 223174
rect -2966 187174 -2346 222618
rect -2966 186618 -2934 187174
rect -2378 186618 -2346 187174
rect -2966 151174 -2346 186618
rect -2966 150618 -2934 151174
rect -2378 150618 -2346 151174
rect -2966 115174 -2346 150618
rect -2966 114618 -2934 115174
rect -2378 114618 -2346 115174
rect -2966 79174 -2346 114618
rect -2966 78618 -2934 79174
rect -2378 78618 -2346 79174
rect -2966 43174 -2346 78618
rect -2966 42618 -2934 43174
rect -2378 42618 -2346 43174
rect -2966 7174 -2346 42618
rect -2966 6618 -2934 7174
rect -2378 6618 -2346 7174
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704282 -1974 704838
rect -1418 704282 -1386 704838
rect -2006 687454 -1386 704282
rect -2006 686898 -1974 687454
rect -1418 686898 -1386 687454
rect -2006 651454 -1386 686898
rect -2006 650898 -1974 651454
rect -1418 650898 -1386 651454
rect -2006 615454 -1386 650898
rect -2006 614898 -1974 615454
rect -1418 614898 -1386 615454
rect -2006 579454 -1386 614898
rect -2006 578898 -1974 579454
rect -1418 578898 -1386 579454
rect -2006 543454 -1386 578898
rect -2006 542898 -1974 543454
rect -1418 542898 -1386 543454
rect -2006 507454 -1386 542898
rect -2006 506898 -1974 507454
rect -1418 506898 -1386 507454
rect -2006 471454 -1386 506898
rect -2006 470898 -1974 471454
rect -1418 470898 -1386 471454
rect -2006 435454 -1386 470898
rect -2006 434898 -1974 435454
rect -1418 434898 -1386 435454
rect -2006 399454 -1386 434898
rect -2006 398898 -1974 399454
rect -1418 398898 -1386 399454
rect -2006 363454 -1386 398898
rect -2006 362898 -1974 363454
rect -1418 362898 -1386 363454
rect -2006 327454 -1386 362898
rect -2006 326898 -1974 327454
rect -1418 326898 -1386 327454
rect -2006 291454 -1386 326898
rect -2006 290898 -1974 291454
rect -1418 290898 -1386 291454
rect -2006 255454 -1386 290898
rect -2006 254898 -1974 255454
rect -1418 254898 -1386 255454
rect -2006 219454 -1386 254898
rect -2006 218898 -1974 219454
rect -1418 218898 -1386 219454
rect -2006 183454 -1386 218898
rect -2006 182898 -1974 183454
rect -1418 182898 -1386 183454
rect -2006 147454 -1386 182898
rect -2006 146898 -1974 147454
rect -1418 146898 -1386 147454
rect -2006 111454 -1386 146898
rect -2006 110898 -1974 111454
rect -1418 110898 -1386 111454
rect -2006 75454 -1386 110898
rect -2006 74898 -1974 75454
rect -1418 74898 -1386 75454
rect -2006 39454 -1386 74898
rect -2006 38898 -1974 39454
rect -1418 38898 -1386 39454
rect -2006 3454 -1386 38898
rect -2006 2898 -1974 3454
rect -1418 2898 -1386 3454
rect -2006 -346 -1386 2898
rect -2006 -902 -1974 -346
rect -1418 -902 -1386 -346
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704282 1826 704838
rect 2382 704282 2414 704838
rect 1794 687454 2414 704282
rect 1794 686898 1826 687454
rect 2382 686898 2414 687454
rect 1794 651454 2414 686898
rect 1794 650898 1826 651454
rect 2382 650898 2414 651454
rect 1794 615454 2414 650898
rect 1794 614898 1826 615454
rect 2382 614898 2414 615454
rect 1794 579454 2414 614898
rect 1794 578898 1826 579454
rect 2382 578898 2414 579454
rect 1794 543454 2414 578898
rect 1794 542898 1826 543454
rect 2382 542898 2414 543454
rect 1794 507454 2414 542898
rect 1794 506898 1826 507454
rect 2382 506898 2414 507454
rect 1794 471454 2414 506898
rect 1794 470898 1826 471454
rect 2382 470898 2414 471454
rect 1794 435454 2414 470898
rect 1794 434898 1826 435454
rect 2382 434898 2414 435454
rect 1794 399454 2414 434898
rect 1794 398898 1826 399454
rect 2382 398898 2414 399454
rect 1794 363454 2414 398898
rect 5514 705798 6134 711590
rect 5514 705242 5546 705798
rect 6102 705242 6134 705798
rect 5514 691174 6134 705242
rect 5514 690618 5546 691174
rect 6102 690618 6134 691174
rect 5514 655174 6134 690618
rect 5514 654618 5546 655174
rect 6102 654618 6134 655174
rect 5514 619174 6134 654618
rect 5514 618618 5546 619174
rect 6102 618618 6134 619174
rect 5514 583174 6134 618618
rect 5514 582618 5546 583174
rect 6102 582618 6134 583174
rect 5514 547174 6134 582618
rect 5514 546618 5546 547174
rect 6102 546618 6134 547174
rect 5514 511174 6134 546618
rect 5514 510618 5546 511174
rect 6102 510618 6134 511174
rect 5514 475174 6134 510618
rect 5514 474618 5546 475174
rect 6102 474618 6134 475174
rect 5514 439174 6134 474618
rect 5514 438618 5546 439174
rect 6102 438618 6134 439174
rect 5514 403174 6134 438618
rect 5514 402618 5546 403174
rect 6102 402618 6134 403174
rect 3739 371380 3805 371381
rect 3739 371316 3740 371380
rect 3804 371316 3805 371380
rect 3739 371315 3805 371316
rect 1794 362898 1826 363454
rect 2382 362898 2414 363454
rect 1794 327454 2414 362898
rect 3555 358460 3621 358461
rect 3555 358396 3556 358460
rect 3620 358396 3621 358460
rect 3555 358395 3621 358396
rect 3371 345404 3437 345405
rect 3371 345340 3372 345404
rect 3436 345340 3437 345404
rect 3371 345339 3437 345340
rect 1794 326898 1826 327454
rect 2382 326898 2414 327454
rect 1794 291454 2414 326898
rect 3374 315893 3434 345339
rect 3558 330309 3618 358395
rect 3742 344725 3802 371315
rect 5514 367174 6134 402618
rect 5514 366618 5546 367174
rect 6102 366618 6134 367174
rect 3739 344724 3805 344725
rect 3739 344660 3740 344724
rect 3804 344660 3805 344724
rect 3739 344659 3805 344660
rect 5514 331174 6134 366618
rect 5514 330618 5546 331174
rect 6102 330618 6134 331174
rect 3555 330308 3621 330309
rect 3555 330244 3556 330308
rect 3620 330244 3621 330308
rect 3555 330243 3621 330244
rect 3739 319292 3805 319293
rect 3739 319228 3740 319292
rect 3804 319228 3805 319292
rect 3739 319227 3805 319228
rect 3371 315892 3437 315893
rect 3371 315828 3372 315892
rect 3436 315828 3437 315892
rect 3371 315827 3437 315828
rect 3555 306236 3621 306237
rect 3555 306172 3556 306236
rect 3620 306172 3621 306236
rect 3555 306171 3621 306172
rect 3371 293180 3437 293181
rect 3371 293116 3372 293180
rect 3436 293116 3437 293180
rect 3371 293115 3437 293116
rect 1794 290898 1826 291454
rect 2382 290898 2414 291454
rect 1794 255454 2414 290898
rect 3374 272645 3434 293115
rect 3558 287061 3618 306171
rect 3742 301477 3802 319227
rect 3739 301476 3805 301477
rect 3739 301412 3740 301476
rect 3804 301412 3805 301476
rect 3739 301411 3805 301412
rect 5514 295174 6134 330618
rect 5514 294618 5546 295174
rect 6102 294618 6134 295174
rect 3555 287060 3621 287061
rect 3555 286996 3556 287060
rect 3620 286996 3621 287060
rect 3555 286995 3621 286996
rect 3371 272644 3437 272645
rect 3371 272580 3372 272644
rect 3436 272580 3437 272644
rect 3371 272579 3437 272580
rect 1794 254898 1826 255454
rect 2382 254898 2414 255454
rect 1794 219454 2414 254898
rect 1794 218898 1826 219454
rect 2382 218898 2414 219454
rect 1794 183454 2414 218898
rect 1794 182898 1826 183454
rect 2382 182898 2414 183454
rect 1794 147454 2414 182898
rect 1794 146898 1826 147454
rect 2382 146898 2414 147454
rect 1794 111454 2414 146898
rect 5514 259174 6134 294618
rect 9234 706758 9854 711590
rect 9234 706202 9266 706758
rect 9822 706202 9854 706758
rect 9234 694894 9854 706202
rect 9234 694338 9266 694894
rect 9822 694338 9854 694894
rect 9234 658894 9854 694338
rect 9234 658338 9266 658894
rect 9822 658338 9854 658894
rect 9234 622894 9854 658338
rect 9234 622338 9266 622894
rect 9822 622338 9854 622894
rect 9234 586894 9854 622338
rect 9234 586338 9266 586894
rect 9822 586338 9854 586894
rect 9234 550894 9854 586338
rect 9234 550338 9266 550894
rect 9822 550338 9854 550894
rect 9234 514894 9854 550338
rect 9234 514338 9266 514894
rect 9822 514338 9854 514894
rect 9234 478894 9854 514338
rect 9234 478338 9266 478894
rect 9822 478338 9854 478894
rect 9234 442894 9854 478338
rect 9234 442338 9266 442894
rect 9822 442338 9854 442894
rect 9234 406894 9854 442338
rect 9234 406338 9266 406894
rect 9822 406338 9854 406894
rect 9234 370894 9854 406338
rect 9234 370338 9266 370894
rect 9822 370338 9854 370894
rect 9234 334894 9854 370338
rect 9234 334338 9266 334894
rect 9822 334338 9854 334894
rect 9234 298894 9854 334338
rect 9234 298338 9266 298894
rect 9822 298338 9854 298894
rect 8155 267204 8221 267205
rect 8155 267140 8156 267204
rect 8220 267140 8221 267204
rect 8155 267139 8221 267140
rect 5514 258618 5546 259174
rect 6102 258618 6134 259174
rect 5514 223174 6134 258618
rect 8158 258229 8218 267139
rect 9234 262894 9854 298338
rect 9234 262338 9266 262894
rect 9822 262338 9854 262894
rect 8155 258228 8221 258229
rect 8155 258164 8156 258228
rect 8220 258164 8221 258228
rect 8155 258163 8221 258164
rect 7419 254148 7485 254149
rect 7419 254084 7420 254148
rect 7484 254084 7485 254148
rect 7419 254083 7485 254084
rect 7422 243813 7482 254083
rect 7419 243812 7485 243813
rect 7419 243748 7420 243812
rect 7484 243748 7485 243812
rect 7419 243747 7485 243748
rect 7419 241092 7485 241093
rect 7419 241028 7420 241092
rect 7484 241028 7485 241092
rect 7419 241027 7485 241028
rect 7422 229397 7482 241027
rect 7419 229396 7485 229397
rect 7419 229332 7420 229396
rect 7484 229332 7485 229396
rect 7419 229331 7485 229332
rect 5514 222618 5546 223174
rect 6102 222618 6134 223174
rect 5514 187174 6134 222618
rect 9234 226894 9854 262338
rect 9234 226338 9266 226894
rect 9822 226338 9854 226894
rect 9234 190894 9854 226338
rect 9234 190338 9266 190894
rect 9822 190338 9854 190894
rect 6315 188868 6381 188869
rect 6315 188804 6316 188868
rect 6380 188804 6381 188868
rect 6315 188803 6381 188804
rect 5514 186618 5546 187174
rect 6102 186618 6134 187174
rect 5514 151174 6134 186618
rect 6318 186149 6378 188803
rect 6315 186148 6381 186149
rect 6315 186084 6316 186148
rect 6380 186084 6381 186148
rect 6315 186083 6381 186084
rect 6315 171732 6381 171733
rect 6315 171668 6316 171732
rect 6380 171668 6381 171732
rect 6315 171667 6381 171668
rect 6318 162893 6378 171667
rect 6315 162892 6381 162893
rect 6315 162828 6316 162892
rect 6380 162828 6381 162892
rect 6315 162827 6381 162828
rect 6315 157316 6381 157317
rect 6315 157252 6316 157316
rect 6380 157252 6381 157316
rect 6315 157251 6381 157252
rect 5514 150618 5546 151174
rect 6102 150618 6134 151174
rect 4843 142900 4909 142901
rect 4843 142836 4844 142900
rect 4908 142836 4909 142900
rect 4843 142835 4909 142836
rect 4846 136781 4906 142835
rect 4843 136780 4909 136781
rect 4843 136716 4844 136780
rect 4908 136716 4909 136780
rect 4843 136715 4909 136716
rect 3371 128484 3437 128485
rect 3371 128420 3372 128484
rect 3436 128420 3437 128484
rect 3371 128419 3437 128420
rect 1794 110898 1826 111454
rect 2382 110898 2414 111454
rect 1794 75454 2414 110898
rect 3374 110669 3434 128419
rect 5514 115174 6134 150618
rect 6318 149837 6378 157251
rect 9234 154894 9854 190338
rect 9234 154338 9266 154894
rect 9822 154338 9854 154894
rect 6315 149836 6381 149837
rect 6315 149772 6316 149836
rect 6380 149772 6381 149836
rect 6315 149771 6381 149772
rect 5514 114618 5546 115174
rect 6102 114618 6134 115174
rect 3555 114068 3621 114069
rect 3555 114004 3556 114068
rect 3620 114004 3621 114068
rect 3555 114003 3621 114004
rect 3371 110668 3437 110669
rect 3371 110604 3372 110668
rect 3436 110604 3437 110668
rect 3371 110603 3437 110604
rect 3558 97613 3618 114003
rect 3555 97612 3621 97613
rect 3555 97548 3556 97612
rect 3620 97548 3621 97612
rect 3555 97547 3621 97548
rect 1794 74898 1826 75454
rect 2382 74898 2414 75454
rect 1794 39454 2414 74898
rect 1794 38898 1826 39454
rect 2382 38898 2414 39454
rect 1794 3454 2414 38898
rect 1794 2898 1826 3454
rect 2382 2898 2414 3454
rect 1794 -346 2414 2898
rect 1794 -902 1826 -346
rect 2382 -902 2414 -346
rect -2966 -1862 -2934 -1306
rect -2378 -1862 -2346 -1306
rect -2966 -1894 -2346 -1862
rect -3926 -2822 -3894 -2266
rect -3338 -2822 -3306 -2266
rect -3926 -2854 -3306 -2822
rect -4886 -3782 -4854 -3226
rect -4298 -3782 -4266 -3226
rect -4886 -3814 -4266 -3782
rect -5846 -4742 -5814 -4186
rect -5258 -4742 -5226 -4186
rect -5846 -4774 -5226 -4742
rect -6806 -5702 -6774 -5146
rect -6218 -5702 -6186 -5146
rect -6806 -5734 -6186 -5702
rect -7766 -6662 -7734 -6106
rect -7178 -6662 -7146 -6106
rect -7766 -6694 -7146 -6662
rect -8726 -7622 -8694 -7066
rect -8138 -7622 -8106 -7066
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 79174 6134 114618
rect 9234 118894 9854 154338
rect 9234 118338 9266 118894
rect 9822 118338 9854 118894
rect 8891 99652 8957 99653
rect 8891 99588 8892 99652
rect 8956 99588 8957 99652
rect 8891 99587 8957 99588
rect 8707 85236 8773 85237
rect 8707 85172 8708 85236
rect 8772 85172 8773 85236
rect 8707 85171 8773 85172
rect 5514 78618 5546 79174
rect 6102 78618 6134 79174
rect 5514 43174 6134 78618
rect 8710 71637 8770 85171
rect 8894 84693 8954 99587
rect 8891 84692 8957 84693
rect 8891 84628 8892 84692
rect 8956 84628 8957 84692
rect 8891 84627 8957 84628
rect 9234 82894 9854 118338
rect 9234 82338 9266 82894
rect 9822 82338 9854 82894
rect 8707 71636 8773 71637
rect 8707 71572 8708 71636
rect 8772 71572 8773 71636
rect 8707 71571 8773 71572
rect 8891 70820 8957 70821
rect 8891 70756 8892 70820
rect 8956 70756 8957 70820
rect 8891 70755 8957 70756
rect 8894 58581 8954 70755
rect 8891 58580 8957 58581
rect 8891 58516 8892 58580
rect 8956 58516 8957 58580
rect 8891 58515 8957 58516
rect 8891 56404 8957 56405
rect 8891 56340 8892 56404
rect 8956 56340 8957 56404
rect 8891 56339 8957 56340
rect 8894 45525 8954 56339
rect 9234 46894 9854 82338
rect 9234 46338 9266 46894
rect 9822 46338 9854 46894
rect 8891 45524 8957 45525
rect 8891 45460 8892 45524
rect 8956 45460 8957 45524
rect 8891 45459 8957 45460
rect 5514 42618 5546 43174
rect 6102 42618 6134 43174
rect 5514 7174 6134 42618
rect 8891 41988 8957 41989
rect 8891 41924 8892 41988
rect 8956 41924 8957 41988
rect 8891 41923 8957 41924
rect 8894 32469 8954 41923
rect 8891 32468 8957 32469
rect 8891 32404 8892 32468
rect 8956 32404 8957 32468
rect 8891 32403 8957 32404
rect 6315 27572 6381 27573
rect 6315 27508 6316 27572
rect 6380 27508 6381 27572
rect 6315 27507 6381 27508
rect 6318 19413 6378 27507
rect 6315 19412 6381 19413
rect 6315 19348 6316 19412
rect 6380 19348 6381 19412
rect 6315 19347 6381 19348
rect 8891 13156 8957 13157
rect 8891 13092 8892 13156
rect 8956 13092 8957 13156
rect 8891 13091 8957 13092
rect 5514 6618 5546 7174
rect 6102 6618 6134 7174
rect 5514 -1306 6134 6618
rect 8894 6493 8954 13091
rect 9234 10894 9854 46338
rect 9234 10338 9266 10894
rect 9822 10338 9854 10894
rect 8891 6492 8957 6493
rect 8891 6428 8892 6492
rect 8956 6428 8957 6492
rect 8891 6427 8957 6428
rect 5514 -1862 5546 -1306
rect 6102 -1862 6134 -1306
rect 5514 -7654 6134 -1862
rect 9234 -2266 9854 10338
rect 9234 -2822 9266 -2266
rect 9822 -2822 9854 -2266
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707162 12986 707718
rect 13542 707162 13574 707718
rect 12954 698614 13574 707162
rect 12954 698058 12986 698614
rect 13542 698058 13574 698614
rect 12954 662614 13574 698058
rect 12954 662058 12986 662614
rect 13542 662058 13574 662614
rect 12954 626614 13574 662058
rect 12954 626058 12986 626614
rect 13542 626058 13574 626614
rect 12954 590614 13574 626058
rect 12954 590058 12986 590614
rect 13542 590058 13574 590614
rect 12954 554614 13574 590058
rect 12954 554058 12986 554614
rect 13542 554058 13574 554614
rect 12954 518614 13574 554058
rect 12954 518058 12986 518614
rect 13542 518058 13574 518614
rect 12954 482614 13574 518058
rect 12954 482058 12986 482614
rect 13542 482058 13574 482614
rect 12954 446614 13574 482058
rect 12954 446058 12986 446614
rect 13542 446058 13574 446614
rect 12954 410614 13574 446058
rect 12954 410058 12986 410614
rect 13542 410058 13574 410614
rect 12954 374614 13574 410058
rect 12954 374058 12986 374614
rect 13542 374058 13574 374614
rect 12954 338614 13574 374058
rect 12954 338058 12986 338614
rect 13542 338058 13574 338614
rect 12954 302614 13574 338058
rect 16674 708678 17294 711590
rect 16674 708122 16706 708678
rect 17262 708122 17294 708678
rect 16674 666334 17294 708122
rect 16674 665778 16706 666334
rect 17262 665778 17294 666334
rect 16674 630334 17294 665778
rect 16674 629778 16706 630334
rect 17262 629778 17294 630334
rect 16674 594334 17294 629778
rect 16674 593778 16706 594334
rect 17262 593778 17294 594334
rect 16674 558334 17294 593778
rect 16674 557778 16706 558334
rect 17262 557778 17294 558334
rect 16674 522334 17294 557778
rect 16674 521778 16706 522334
rect 17262 521778 17294 522334
rect 16674 486334 17294 521778
rect 16674 485778 16706 486334
rect 17262 485778 17294 486334
rect 16674 450334 17294 485778
rect 16674 449778 16706 450334
rect 17262 449778 17294 450334
rect 16674 414334 17294 449778
rect 16674 413778 16706 414334
rect 17262 413778 17294 414334
rect 16674 378334 17294 413778
rect 16674 377778 16706 378334
rect 17262 377778 17294 378334
rect 16674 342334 17294 377778
rect 16674 341778 16706 342334
rect 17262 341778 17294 342334
rect 16208 327454 16528 327486
rect 16208 327218 16250 327454
rect 16486 327218 16528 327454
rect 16208 327134 16528 327218
rect 16208 326898 16250 327134
rect 16486 326898 16528 327134
rect 16208 326866 16528 326898
rect 12954 302058 12986 302614
rect 13542 302058 13574 302614
rect 12954 266614 13574 302058
rect 16674 306334 17294 341778
rect 16674 305778 16706 306334
rect 17262 305778 17294 306334
rect 16208 291454 16528 291486
rect 16208 291218 16250 291454
rect 16486 291218 16528 291454
rect 16208 291134 16528 291218
rect 16208 290898 16250 291134
rect 16486 290898 16528 291134
rect 16208 290866 16528 290898
rect 12954 266058 12986 266614
rect 13542 266058 13574 266614
rect 12954 230614 13574 266058
rect 16674 270334 17294 305778
rect 16674 269778 16706 270334
rect 17262 269778 17294 270334
rect 16208 255454 16528 255486
rect 16208 255218 16250 255454
rect 16486 255218 16528 255454
rect 16208 255134 16528 255218
rect 16208 254898 16250 255134
rect 16486 254898 16528 255134
rect 16208 254866 16528 254898
rect 12954 230058 12986 230614
rect 13542 230058 13574 230614
rect 12954 194614 13574 230058
rect 16674 234334 17294 269778
rect 16674 233778 16706 234334
rect 17262 233778 17294 234334
rect 16208 219454 16528 219486
rect 16208 219218 16250 219454
rect 16486 219218 16528 219454
rect 16208 219134 16528 219218
rect 16208 218898 16250 219134
rect 16486 218898 16528 219134
rect 16208 218866 16528 218898
rect 12954 194058 12986 194614
rect 13542 194058 13574 194614
rect 12954 158614 13574 194058
rect 16674 198334 17294 233778
rect 16674 197778 16706 198334
rect 17262 197778 17294 198334
rect 16208 183454 16528 183486
rect 16208 183218 16250 183454
rect 16486 183218 16528 183454
rect 16208 183134 16528 183218
rect 16208 182898 16250 183134
rect 16486 182898 16528 183134
rect 16208 182866 16528 182898
rect 12954 158058 12986 158614
rect 13542 158058 13574 158614
rect 12954 122614 13574 158058
rect 16674 162334 17294 197778
rect 16674 161778 16706 162334
rect 17262 161778 17294 162334
rect 16208 147454 16528 147486
rect 16208 147218 16250 147454
rect 16486 147218 16528 147454
rect 16208 147134 16528 147218
rect 16208 146898 16250 147134
rect 16486 146898 16528 147134
rect 16208 146866 16528 146898
rect 12954 122058 12986 122614
rect 13542 122058 13574 122614
rect 12954 86614 13574 122058
rect 16674 126334 17294 161778
rect 16674 125778 16706 126334
rect 17262 125778 17294 126334
rect 16208 111454 16528 111486
rect 16208 111218 16250 111454
rect 16486 111218 16528 111454
rect 16208 111134 16528 111218
rect 16208 110898 16250 111134
rect 16486 110898 16528 111134
rect 16208 110866 16528 110898
rect 12954 86058 12986 86614
rect 13542 86058 13574 86614
rect 12954 50614 13574 86058
rect 16674 90334 17294 125778
rect 16674 89778 16706 90334
rect 17262 89778 17294 90334
rect 16208 75454 16528 75486
rect 16208 75218 16250 75454
rect 16486 75218 16528 75454
rect 16208 75134 16528 75218
rect 16208 74898 16250 75134
rect 16486 74898 16528 75134
rect 16208 74866 16528 74898
rect 12954 50058 12986 50614
rect 13542 50058 13574 50614
rect 12954 14614 13574 50058
rect 16674 54334 17294 89778
rect 16674 53778 16706 54334
rect 17262 53778 17294 54334
rect 16208 39454 16528 39486
rect 16208 39218 16250 39454
rect 16486 39218 16528 39454
rect 16208 39134 16528 39218
rect 16208 38898 16250 39134
rect 16486 38898 16528 39134
rect 16208 38866 16528 38898
rect 12954 14058 12986 14614
rect 13542 14058 13574 14614
rect 12954 -3226 13574 14058
rect 12954 -3782 12986 -3226
rect 13542 -3782 13574 -3226
rect 12954 -7654 13574 -3782
rect 16674 18334 17294 53778
rect 16674 17778 16706 18334
rect 17262 17778 17294 18334
rect 16674 -4186 17294 17778
rect 16674 -4742 16706 -4186
rect 17262 -4742 17294 -4186
rect 16674 -7654 17294 -4742
rect 20394 709638 21014 711590
rect 20394 709082 20426 709638
rect 20982 709082 21014 709638
rect 20394 670054 21014 709082
rect 20394 669498 20426 670054
rect 20982 669498 21014 670054
rect 20394 634054 21014 669498
rect 20394 633498 20426 634054
rect 20982 633498 21014 634054
rect 20394 598054 21014 633498
rect 20394 597498 20426 598054
rect 20982 597498 21014 598054
rect 20394 562054 21014 597498
rect 20394 561498 20426 562054
rect 20982 561498 21014 562054
rect 20394 526054 21014 561498
rect 20394 525498 20426 526054
rect 20982 525498 21014 526054
rect 20394 490054 21014 525498
rect 20394 489498 20426 490054
rect 20982 489498 21014 490054
rect 20394 454054 21014 489498
rect 20394 453498 20426 454054
rect 20982 453498 21014 454054
rect 20394 418054 21014 453498
rect 20394 417498 20426 418054
rect 20982 417498 21014 418054
rect 20394 382054 21014 417498
rect 20394 381498 20426 382054
rect 20982 381498 21014 382054
rect 20394 346054 21014 381498
rect 20394 345498 20426 346054
rect 20982 345498 21014 346054
rect 20394 310054 21014 345498
rect 20394 309498 20426 310054
rect 20982 309498 21014 310054
rect 20394 274054 21014 309498
rect 20394 273498 20426 274054
rect 20982 273498 21014 274054
rect 20394 238054 21014 273498
rect 20394 237498 20426 238054
rect 20982 237498 21014 238054
rect 20394 202054 21014 237498
rect 20394 201498 20426 202054
rect 20982 201498 21014 202054
rect 20394 166054 21014 201498
rect 20394 165498 20426 166054
rect 20982 165498 21014 166054
rect 20394 130054 21014 165498
rect 20394 129498 20426 130054
rect 20982 129498 21014 130054
rect 20394 94054 21014 129498
rect 20394 93498 20426 94054
rect 20982 93498 21014 94054
rect 20394 58054 21014 93498
rect 20394 57498 20426 58054
rect 20982 57498 21014 58054
rect 20394 22054 21014 57498
rect 20394 21498 20426 22054
rect 20982 21498 21014 22054
rect 20394 -5146 21014 21498
rect 20394 -5702 20426 -5146
rect 20982 -5702 21014 -5146
rect 20394 -7654 21014 -5702
rect 24114 710598 24734 711590
rect 24114 710042 24146 710598
rect 24702 710042 24734 710598
rect 24114 673774 24734 710042
rect 24114 673218 24146 673774
rect 24702 673218 24734 673774
rect 24114 637774 24734 673218
rect 24114 637218 24146 637774
rect 24702 637218 24734 637774
rect 24114 601774 24734 637218
rect 24114 601218 24146 601774
rect 24702 601218 24734 601774
rect 24114 565774 24734 601218
rect 24114 565218 24146 565774
rect 24702 565218 24734 565774
rect 24114 529774 24734 565218
rect 24114 529218 24146 529774
rect 24702 529218 24734 529774
rect 24114 493774 24734 529218
rect 24114 493218 24146 493774
rect 24702 493218 24734 493774
rect 24114 457774 24734 493218
rect 24114 457218 24146 457774
rect 24702 457218 24734 457774
rect 24114 421774 24734 457218
rect 24114 421218 24146 421774
rect 24702 421218 24734 421774
rect 24114 385774 24734 421218
rect 24114 385218 24146 385774
rect 24702 385218 24734 385774
rect 24114 349774 24734 385218
rect 24114 349218 24146 349774
rect 24702 349218 24734 349774
rect 24114 313774 24734 349218
rect 24114 313218 24146 313774
rect 24702 313218 24734 313774
rect 24114 277774 24734 313218
rect 24114 277218 24146 277774
rect 24702 277218 24734 277774
rect 24114 241774 24734 277218
rect 24114 241218 24146 241774
rect 24702 241218 24734 241774
rect 24114 205774 24734 241218
rect 24114 205218 24146 205774
rect 24702 205218 24734 205774
rect 24114 169774 24734 205218
rect 24114 169218 24146 169774
rect 24702 169218 24734 169774
rect 24114 133774 24734 169218
rect 24114 133218 24146 133774
rect 24702 133218 24734 133774
rect 24114 97774 24734 133218
rect 24114 97218 24146 97774
rect 24702 97218 24734 97774
rect 24114 61774 24734 97218
rect 24114 61218 24146 61774
rect 24702 61218 24734 61774
rect 24114 25774 24734 61218
rect 24114 25218 24146 25774
rect 24702 25218 24734 25774
rect 24114 -6106 24734 25218
rect 24114 -6662 24146 -6106
rect 24702 -6662 24734 -6106
rect 24114 -7654 24734 -6662
rect 27834 711558 28454 711590
rect 27834 711002 27866 711558
rect 28422 711002 28454 711558
rect 27834 677494 28454 711002
rect 27834 676938 27866 677494
rect 28422 676938 28454 677494
rect 27834 641494 28454 676938
rect 27834 640938 27866 641494
rect 28422 640938 28454 641494
rect 27834 605494 28454 640938
rect 27834 604938 27866 605494
rect 28422 604938 28454 605494
rect 27834 569494 28454 604938
rect 27834 568938 27866 569494
rect 28422 568938 28454 569494
rect 27834 533494 28454 568938
rect 27834 532938 27866 533494
rect 28422 532938 28454 533494
rect 27834 497494 28454 532938
rect 27834 496938 27866 497494
rect 28422 496938 28454 497494
rect 27834 461494 28454 496938
rect 27834 460938 27866 461494
rect 28422 460938 28454 461494
rect 27834 425494 28454 460938
rect 27834 424938 27866 425494
rect 28422 424938 28454 425494
rect 27834 389494 28454 424938
rect 27834 388938 27866 389494
rect 28422 388938 28454 389494
rect 27834 353494 28454 388938
rect 27834 352938 27866 353494
rect 28422 352938 28454 353494
rect 27834 317494 28454 352938
rect 37794 704838 38414 711590
rect 37794 704282 37826 704838
rect 38382 704282 38414 704838
rect 37794 687454 38414 704282
rect 37794 686898 37826 687454
rect 38382 686898 38414 687454
rect 37794 651454 38414 686898
rect 37794 650898 37826 651454
rect 38382 650898 38414 651454
rect 37794 615454 38414 650898
rect 37794 614898 37826 615454
rect 38382 614898 38414 615454
rect 37794 579454 38414 614898
rect 37794 578898 37826 579454
rect 38382 578898 38414 579454
rect 37794 543454 38414 578898
rect 37794 542898 37826 543454
rect 38382 542898 38414 543454
rect 37794 507454 38414 542898
rect 37794 506898 37826 507454
rect 38382 506898 38414 507454
rect 37794 471454 38414 506898
rect 37794 470898 37826 471454
rect 38382 470898 38414 471454
rect 37794 435454 38414 470898
rect 37794 434898 37826 435454
rect 38382 434898 38414 435454
rect 37794 399454 38414 434898
rect 37794 398898 37826 399454
rect 38382 398898 38414 399454
rect 37794 363454 38414 398898
rect 37794 362898 37826 363454
rect 38382 362898 38414 363454
rect 31568 331174 31888 331206
rect 31568 330938 31610 331174
rect 31846 330938 31888 331174
rect 31568 330854 31888 330938
rect 31568 330618 31610 330854
rect 31846 330618 31888 330854
rect 31568 330586 31888 330618
rect 27834 316938 27866 317494
rect 28422 316938 28454 317494
rect 27834 281494 28454 316938
rect 37794 327454 38414 362898
rect 37794 326898 37826 327454
rect 38382 326898 38414 327454
rect 31568 295174 31888 295206
rect 31568 294938 31610 295174
rect 31846 294938 31888 295174
rect 31568 294854 31888 294938
rect 31568 294618 31610 294854
rect 31846 294618 31888 294854
rect 31568 294586 31888 294618
rect 27834 280938 27866 281494
rect 28422 280938 28454 281494
rect 27834 245494 28454 280938
rect 37794 291454 38414 326898
rect 37794 290898 37826 291454
rect 38382 290898 38414 291454
rect 31568 259174 31888 259206
rect 31568 258938 31610 259174
rect 31846 258938 31888 259174
rect 31568 258854 31888 258938
rect 31568 258618 31610 258854
rect 31846 258618 31888 258854
rect 31568 258586 31888 258618
rect 27834 244938 27866 245494
rect 28422 244938 28454 245494
rect 27834 209494 28454 244938
rect 37794 255454 38414 290898
rect 37794 254898 37826 255454
rect 38382 254898 38414 255454
rect 31568 223174 31888 223206
rect 31568 222938 31610 223174
rect 31846 222938 31888 223174
rect 31568 222854 31888 222938
rect 31568 222618 31610 222854
rect 31846 222618 31888 222854
rect 31568 222586 31888 222618
rect 27834 208938 27866 209494
rect 28422 208938 28454 209494
rect 27834 173494 28454 208938
rect 37794 219454 38414 254898
rect 37794 218898 37826 219454
rect 38382 218898 38414 219454
rect 31568 187174 31888 187206
rect 31568 186938 31610 187174
rect 31846 186938 31888 187174
rect 31568 186854 31888 186938
rect 31568 186618 31610 186854
rect 31846 186618 31888 186854
rect 31568 186586 31888 186618
rect 27834 172938 27866 173494
rect 28422 172938 28454 173494
rect 27834 137494 28454 172938
rect 37794 183454 38414 218898
rect 37794 182898 37826 183454
rect 38382 182898 38414 183454
rect 31568 151174 31888 151206
rect 31568 150938 31610 151174
rect 31846 150938 31888 151174
rect 31568 150854 31888 150938
rect 31568 150618 31610 150854
rect 31846 150618 31888 150854
rect 31568 150586 31888 150618
rect 27834 136938 27866 137494
rect 28422 136938 28454 137494
rect 27834 101494 28454 136938
rect 37794 147454 38414 182898
rect 37794 146898 37826 147454
rect 38382 146898 38414 147454
rect 31568 115174 31888 115206
rect 31568 114938 31610 115174
rect 31846 114938 31888 115174
rect 31568 114854 31888 114938
rect 31568 114618 31610 114854
rect 31846 114618 31888 114854
rect 31568 114586 31888 114618
rect 27834 100938 27866 101494
rect 28422 100938 28454 101494
rect 27834 65494 28454 100938
rect 37794 111454 38414 146898
rect 37794 110898 37826 111454
rect 38382 110898 38414 111454
rect 31568 79174 31888 79206
rect 31568 78938 31610 79174
rect 31846 78938 31888 79174
rect 31568 78854 31888 78938
rect 31568 78618 31610 78854
rect 31846 78618 31888 78854
rect 31568 78586 31888 78618
rect 27834 64938 27866 65494
rect 28422 64938 28454 65494
rect 27834 29494 28454 64938
rect 37794 75454 38414 110898
rect 37794 74898 37826 75454
rect 38382 74898 38414 75454
rect 31568 43174 31888 43206
rect 31568 42938 31610 43174
rect 31846 42938 31888 43174
rect 31568 42854 31888 42938
rect 31568 42618 31610 42854
rect 31846 42618 31888 42854
rect 31568 42586 31888 42618
rect 27834 28938 27866 29494
rect 28422 28938 28454 29494
rect 27834 -7066 28454 28938
rect 37794 39454 38414 74898
rect 37794 38898 37826 39454
rect 38382 38898 38414 39454
rect 31568 7174 31888 7206
rect 31568 6938 31610 7174
rect 31846 6938 31888 7174
rect 31568 6854 31888 6938
rect 31568 6618 31610 6854
rect 31846 6618 31888 6854
rect 31568 6586 31888 6618
rect 37794 3454 38414 38898
rect 34835 3228 34901 3229
rect 34835 3164 34836 3228
rect 34900 3164 34901 3228
rect 34835 3163 34901 3164
rect 34838 2549 34898 3163
rect 37794 2898 37826 3454
rect 38382 2898 38414 3454
rect 34835 2548 34901 2549
rect 34835 2484 34836 2548
rect 34900 2484 34901 2548
rect 34835 2483 34901 2484
rect 27834 -7622 27866 -7066
rect 28422 -7622 28454 -7066
rect 27834 -7654 28454 -7622
rect 37794 -346 38414 2898
rect 37794 -902 37826 -346
rect 38382 -902 38414 -346
rect 37794 -7654 38414 -902
rect 41514 705798 42134 711590
rect 41514 705242 41546 705798
rect 42102 705242 42134 705798
rect 41514 691174 42134 705242
rect 41514 690618 41546 691174
rect 42102 690618 42134 691174
rect 41514 655174 42134 690618
rect 41514 654618 41546 655174
rect 42102 654618 42134 655174
rect 41514 619174 42134 654618
rect 41514 618618 41546 619174
rect 42102 618618 42134 619174
rect 41514 583174 42134 618618
rect 41514 582618 41546 583174
rect 42102 582618 42134 583174
rect 41514 547174 42134 582618
rect 41514 546618 41546 547174
rect 42102 546618 42134 547174
rect 41514 511174 42134 546618
rect 41514 510618 41546 511174
rect 42102 510618 42134 511174
rect 41514 475174 42134 510618
rect 41514 474618 41546 475174
rect 42102 474618 42134 475174
rect 41514 439174 42134 474618
rect 41514 438618 41546 439174
rect 42102 438618 42134 439174
rect 41514 403174 42134 438618
rect 41514 402618 41546 403174
rect 42102 402618 42134 403174
rect 41514 367174 42134 402618
rect 41514 366618 41546 367174
rect 42102 366618 42134 367174
rect 41514 331174 42134 366618
rect 41514 330618 41546 331174
rect 42102 330618 42134 331174
rect 41514 295174 42134 330618
rect 41514 294618 41546 295174
rect 42102 294618 42134 295174
rect 41514 259174 42134 294618
rect 41514 258618 41546 259174
rect 42102 258618 42134 259174
rect 41514 223174 42134 258618
rect 41514 222618 41546 223174
rect 42102 222618 42134 223174
rect 41514 187174 42134 222618
rect 41514 186618 41546 187174
rect 42102 186618 42134 187174
rect 41514 151174 42134 186618
rect 41514 150618 41546 151174
rect 42102 150618 42134 151174
rect 41514 115174 42134 150618
rect 41514 114618 41546 115174
rect 42102 114618 42134 115174
rect 41514 79174 42134 114618
rect 41514 78618 41546 79174
rect 42102 78618 42134 79174
rect 41514 43174 42134 78618
rect 41514 42618 41546 43174
rect 42102 42618 42134 43174
rect 41514 7174 42134 42618
rect 41514 6618 41546 7174
rect 42102 6618 42134 7174
rect 41514 -1306 42134 6618
rect 41514 -1862 41546 -1306
rect 42102 -1862 42134 -1306
rect 41514 -7654 42134 -1862
rect 45234 706758 45854 711590
rect 45234 706202 45266 706758
rect 45822 706202 45854 706758
rect 45234 694894 45854 706202
rect 45234 694338 45266 694894
rect 45822 694338 45854 694894
rect 45234 658894 45854 694338
rect 45234 658338 45266 658894
rect 45822 658338 45854 658894
rect 45234 622894 45854 658338
rect 45234 622338 45266 622894
rect 45822 622338 45854 622894
rect 45234 586894 45854 622338
rect 45234 586338 45266 586894
rect 45822 586338 45854 586894
rect 45234 550894 45854 586338
rect 45234 550338 45266 550894
rect 45822 550338 45854 550894
rect 45234 514894 45854 550338
rect 45234 514338 45266 514894
rect 45822 514338 45854 514894
rect 45234 478894 45854 514338
rect 45234 478338 45266 478894
rect 45822 478338 45854 478894
rect 45234 442894 45854 478338
rect 45234 442338 45266 442894
rect 45822 442338 45854 442894
rect 45234 406894 45854 442338
rect 45234 406338 45266 406894
rect 45822 406338 45854 406894
rect 45234 370894 45854 406338
rect 45234 370338 45266 370894
rect 45822 370338 45854 370894
rect 45234 334894 45854 370338
rect 45234 334338 45266 334894
rect 45822 334338 45854 334894
rect 45234 298894 45854 334338
rect 48954 707718 49574 711590
rect 48954 707162 48986 707718
rect 49542 707162 49574 707718
rect 48954 698614 49574 707162
rect 48954 698058 48986 698614
rect 49542 698058 49574 698614
rect 48954 662614 49574 698058
rect 48954 662058 48986 662614
rect 49542 662058 49574 662614
rect 48954 626614 49574 662058
rect 48954 626058 48986 626614
rect 49542 626058 49574 626614
rect 48954 590614 49574 626058
rect 48954 590058 48986 590614
rect 49542 590058 49574 590614
rect 48954 554614 49574 590058
rect 48954 554058 48986 554614
rect 49542 554058 49574 554614
rect 48954 518614 49574 554058
rect 48954 518058 48986 518614
rect 49542 518058 49574 518614
rect 48954 482614 49574 518058
rect 48954 482058 48986 482614
rect 49542 482058 49574 482614
rect 48954 446614 49574 482058
rect 48954 446058 48986 446614
rect 49542 446058 49574 446614
rect 48954 410614 49574 446058
rect 48954 410058 48986 410614
rect 49542 410058 49574 410614
rect 48954 374614 49574 410058
rect 48954 374058 48986 374614
rect 49542 374058 49574 374614
rect 48954 338614 49574 374058
rect 48954 338058 48986 338614
rect 49542 338058 49574 338614
rect 46928 327454 47248 327486
rect 46928 327218 46970 327454
rect 47206 327218 47248 327454
rect 46928 327134 47248 327218
rect 46928 326898 46970 327134
rect 47206 326898 47248 327134
rect 46928 326866 47248 326898
rect 45234 298338 45266 298894
rect 45822 298338 45854 298894
rect 45234 262894 45854 298338
rect 48954 302614 49574 338058
rect 48954 302058 48986 302614
rect 49542 302058 49574 302614
rect 46928 291454 47248 291486
rect 46928 291218 46970 291454
rect 47206 291218 47248 291454
rect 46928 291134 47248 291218
rect 46928 290898 46970 291134
rect 47206 290898 47248 291134
rect 46928 290866 47248 290898
rect 45234 262338 45266 262894
rect 45822 262338 45854 262894
rect 45234 226894 45854 262338
rect 48954 266614 49574 302058
rect 48954 266058 48986 266614
rect 49542 266058 49574 266614
rect 46928 255454 47248 255486
rect 46928 255218 46970 255454
rect 47206 255218 47248 255454
rect 46928 255134 47248 255218
rect 46928 254898 46970 255134
rect 47206 254898 47248 255134
rect 46928 254866 47248 254898
rect 45234 226338 45266 226894
rect 45822 226338 45854 226894
rect 45234 190894 45854 226338
rect 48954 230614 49574 266058
rect 48954 230058 48986 230614
rect 49542 230058 49574 230614
rect 46928 219454 47248 219486
rect 46928 219218 46970 219454
rect 47206 219218 47248 219454
rect 46928 219134 47248 219218
rect 46928 218898 46970 219134
rect 47206 218898 47248 219134
rect 46928 218866 47248 218898
rect 45234 190338 45266 190894
rect 45822 190338 45854 190894
rect 45234 154894 45854 190338
rect 48954 194614 49574 230058
rect 48954 194058 48986 194614
rect 49542 194058 49574 194614
rect 46928 183454 47248 183486
rect 46928 183218 46970 183454
rect 47206 183218 47248 183454
rect 46928 183134 47248 183218
rect 46928 182898 46970 183134
rect 47206 182898 47248 183134
rect 46928 182866 47248 182898
rect 45234 154338 45266 154894
rect 45822 154338 45854 154894
rect 45234 118894 45854 154338
rect 48954 158614 49574 194058
rect 48954 158058 48986 158614
rect 49542 158058 49574 158614
rect 46928 147454 47248 147486
rect 46928 147218 46970 147454
rect 47206 147218 47248 147454
rect 46928 147134 47248 147218
rect 46928 146898 46970 147134
rect 47206 146898 47248 147134
rect 46928 146866 47248 146898
rect 45234 118338 45266 118894
rect 45822 118338 45854 118894
rect 45234 82894 45854 118338
rect 48954 122614 49574 158058
rect 48954 122058 48986 122614
rect 49542 122058 49574 122614
rect 46928 111454 47248 111486
rect 46928 111218 46970 111454
rect 47206 111218 47248 111454
rect 46928 111134 47248 111218
rect 46928 110898 46970 111134
rect 47206 110898 47248 111134
rect 46928 110866 47248 110898
rect 45234 82338 45266 82894
rect 45822 82338 45854 82894
rect 45234 46894 45854 82338
rect 48954 86614 49574 122058
rect 48954 86058 48986 86614
rect 49542 86058 49574 86614
rect 46928 75454 47248 75486
rect 46928 75218 46970 75454
rect 47206 75218 47248 75454
rect 46928 75134 47248 75218
rect 46928 74898 46970 75134
rect 47206 74898 47248 75134
rect 46928 74866 47248 74898
rect 45234 46338 45266 46894
rect 45822 46338 45854 46894
rect 45234 10894 45854 46338
rect 48954 50614 49574 86058
rect 48954 50058 48986 50614
rect 49542 50058 49574 50614
rect 46928 39454 47248 39486
rect 46928 39218 46970 39454
rect 47206 39218 47248 39454
rect 46928 39134 47248 39218
rect 46928 38898 46970 39134
rect 47206 38898 47248 39134
rect 46928 38866 47248 38898
rect 45234 10338 45266 10894
rect 45822 10338 45854 10894
rect 45234 -2266 45854 10338
rect 48954 14614 49574 50058
rect 48954 14058 48986 14614
rect 49542 14058 49574 14614
rect 47899 3908 47965 3909
rect 47899 3844 47900 3908
rect 47964 3844 47965 3908
rect 47899 3843 47965 3844
rect 47902 2685 47962 3843
rect 47899 2684 47965 2685
rect 47899 2620 47900 2684
rect 47964 2620 47965 2684
rect 47899 2619 47965 2620
rect 45234 -2822 45266 -2266
rect 45822 -2822 45854 -2266
rect 45234 -7654 45854 -2822
rect 48954 -3226 49574 14058
rect 48954 -3782 48986 -3226
rect 49542 -3782 49574 -3226
rect 48954 -7654 49574 -3782
rect 52674 708678 53294 711590
rect 52674 708122 52706 708678
rect 53262 708122 53294 708678
rect 52674 666334 53294 708122
rect 52674 665778 52706 666334
rect 53262 665778 53294 666334
rect 52674 630334 53294 665778
rect 52674 629778 52706 630334
rect 53262 629778 53294 630334
rect 52674 594334 53294 629778
rect 52674 593778 52706 594334
rect 53262 593778 53294 594334
rect 52674 558334 53294 593778
rect 52674 557778 52706 558334
rect 53262 557778 53294 558334
rect 52674 522334 53294 557778
rect 52674 521778 52706 522334
rect 53262 521778 53294 522334
rect 52674 486334 53294 521778
rect 52674 485778 52706 486334
rect 53262 485778 53294 486334
rect 52674 450334 53294 485778
rect 52674 449778 52706 450334
rect 53262 449778 53294 450334
rect 52674 414334 53294 449778
rect 52674 413778 52706 414334
rect 53262 413778 53294 414334
rect 52674 378334 53294 413778
rect 52674 377778 52706 378334
rect 53262 377778 53294 378334
rect 52674 342334 53294 377778
rect 52674 341778 52706 342334
rect 53262 341778 53294 342334
rect 52674 306334 53294 341778
rect 52674 305778 52706 306334
rect 53262 305778 53294 306334
rect 52674 270334 53294 305778
rect 52674 269778 52706 270334
rect 53262 269778 53294 270334
rect 52674 234334 53294 269778
rect 52674 233778 52706 234334
rect 53262 233778 53294 234334
rect 52674 198334 53294 233778
rect 52674 197778 52706 198334
rect 53262 197778 53294 198334
rect 52674 162334 53294 197778
rect 52674 161778 52706 162334
rect 53262 161778 53294 162334
rect 52674 126334 53294 161778
rect 52674 125778 52706 126334
rect 53262 125778 53294 126334
rect 52674 90334 53294 125778
rect 52674 89778 52706 90334
rect 53262 89778 53294 90334
rect 52674 54334 53294 89778
rect 52674 53778 52706 54334
rect 53262 53778 53294 54334
rect 52674 18334 53294 53778
rect 52674 17778 52706 18334
rect 53262 17778 53294 18334
rect 52674 -4186 53294 17778
rect 52674 -4742 52706 -4186
rect 53262 -4742 53294 -4186
rect 52674 -7654 53294 -4742
rect 56394 709638 57014 711590
rect 56394 709082 56426 709638
rect 56982 709082 57014 709638
rect 56394 670054 57014 709082
rect 56394 669498 56426 670054
rect 56982 669498 57014 670054
rect 56394 634054 57014 669498
rect 56394 633498 56426 634054
rect 56982 633498 57014 634054
rect 56394 598054 57014 633498
rect 56394 597498 56426 598054
rect 56982 597498 57014 598054
rect 56394 562054 57014 597498
rect 56394 561498 56426 562054
rect 56982 561498 57014 562054
rect 56394 526054 57014 561498
rect 56394 525498 56426 526054
rect 56982 525498 57014 526054
rect 56394 490054 57014 525498
rect 56394 489498 56426 490054
rect 56982 489498 57014 490054
rect 56394 454054 57014 489498
rect 56394 453498 56426 454054
rect 56982 453498 57014 454054
rect 56394 418054 57014 453498
rect 56394 417498 56426 418054
rect 56982 417498 57014 418054
rect 56394 382054 57014 417498
rect 56394 381498 56426 382054
rect 56982 381498 57014 382054
rect 56394 346054 57014 381498
rect 56394 345498 56426 346054
rect 56982 345498 57014 346054
rect 56394 310054 57014 345498
rect 56394 309498 56426 310054
rect 56982 309498 57014 310054
rect 56394 274054 57014 309498
rect 56394 273498 56426 274054
rect 56982 273498 57014 274054
rect 56394 238054 57014 273498
rect 56394 237498 56426 238054
rect 56982 237498 57014 238054
rect 56394 202054 57014 237498
rect 56394 201498 56426 202054
rect 56982 201498 57014 202054
rect 56394 166054 57014 201498
rect 56394 165498 56426 166054
rect 56982 165498 57014 166054
rect 56394 130054 57014 165498
rect 56394 129498 56426 130054
rect 56982 129498 57014 130054
rect 56394 94054 57014 129498
rect 56394 93498 56426 94054
rect 56982 93498 57014 94054
rect 56394 58054 57014 93498
rect 56394 57498 56426 58054
rect 56982 57498 57014 58054
rect 56394 22054 57014 57498
rect 56394 21498 56426 22054
rect 56982 21498 57014 22054
rect 56394 -5146 57014 21498
rect 60114 710598 60734 711590
rect 60114 710042 60146 710598
rect 60702 710042 60734 710598
rect 60114 673774 60734 710042
rect 60114 673218 60146 673774
rect 60702 673218 60734 673774
rect 60114 637774 60734 673218
rect 60114 637218 60146 637774
rect 60702 637218 60734 637774
rect 60114 601774 60734 637218
rect 60114 601218 60146 601774
rect 60702 601218 60734 601774
rect 60114 565774 60734 601218
rect 60114 565218 60146 565774
rect 60702 565218 60734 565774
rect 60114 529774 60734 565218
rect 60114 529218 60146 529774
rect 60702 529218 60734 529774
rect 60114 493774 60734 529218
rect 60114 493218 60146 493774
rect 60702 493218 60734 493774
rect 60114 457774 60734 493218
rect 60114 457218 60146 457774
rect 60702 457218 60734 457774
rect 60114 421774 60734 457218
rect 60114 421218 60146 421774
rect 60702 421218 60734 421774
rect 60114 385774 60734 421218
rect 60114 385218 60146 385774
rect 60702 385218 60734 385774
rect 60114 349774 60734 385218
rect 60114 349218 60146 349774
rect 60702 349218 60734 349774
rect 60114 313774 60734 349218
rect 63834 711558 64454 711590
rect 63834 711002 63866 711558
rect 64422 711002 64454 711558
rect 63834 677494 64454 711002
rect 63834 676938 63866 677494
rect 64422 676938 64454 677494
rect 63834 641494 64454 676938
rect 63834 640938 63866 641494
rect 64422 640938 64454 641494
rect 63834 605494 64454 640938
rect 63834 604938 63866 605494
rect 64422 604938 64454 605494
rect 63834 569494 64454 604938
rect 63834 568938 63866 569494
rect 64422 568938 64454 569494
rect 63834 533494 64454 568938
rect 63834 532938 63866 533494
rect 64422 532938 64454 533494
rect 63834 497494 64454 532938
rect 63834 496938 63866 497494
rect 64422 496938 64454 497494
rect 63834 461494 64454 496938
rect 63834 460938 63866 461494
rect 64422 460938 64454 461494
rect 63834 425494 64454 460938
rect 63834 424938 63866 425494
rect 64422 424938 64454 425494
rect 63834 389494 64454 424938
rect 63834 388938 63866 389494
rect 64422 388938 64454 389494
rect 63834 353494 64454 388938
rect 63834 352938 63866 353494
rect 64422 352938 64454 353494
rect 62288 331174 62608 331206
rect 62288 330938 62330 331174
rect 62566 330938 62608 331174
rect 62288 330854 62608 330938
rect 62288 330618 62330 330854
rect 62566 330618 62608 330854
rect 62288 330586 62608 330618
rect 60114 313218 60146 313774
rect 60702 313218 60734 313774
rect 60114 277774 60734 313218
rect 63834 317494 64454 352938
rect 63834 316938 63866 317494
rect 64422 316938 64454 317494
rect 62288 295174 62608 295206
rect 62288 294938 62330 295174
rect 62566 294938 62608 295174
rect 62288 294854 62608 294938
rect 62288 294618 62330 294854
rect 62566 294618 62608 294854
rect 62288 294586 62608 294618
rect 60114 277218 60146 277774
rect 60702 277218 60734 277774
rect 60114 241774 60734 277218
rect 63834 281494 64454 316938
rect 63834 280938 63866 281494
rect 64422 280938 64454 281494
rect 62288 259174 62608 259206
rect 62288 258938 62330 259174
rect 62566 258938 62608 259174
rect 62288 258854 62608 258938
rect 62288 258618 62330 258854
rect 62566 258618 62608 258854
rect 62288 258586 62608 258618
rect 60114 241218 60146 241774
rect 60702 241218 60734 241774
rect 60114 205774 60734 241218
rect 63834 245494 64454 280938
rect 63834 244938 63866 245494
rect 64422 244938 64454 245494
rect 62288 223174 62608 223206
rect 62288 222938 62330 223174
rect 62566 222938 62608 223174
rect 62288 222854 62608 222938
rect 62288 222618 62330 222854
rect 62566 222618 62608 222854
rect 62288 222586 62608 222618
rect 60114 205218 60146 205774
rect 60702 205218 60734 205774
rect 60114 169774 60734 205218
rect 63834 209494 64454 244938
rect 63834 208938 63866 209494
rect 64422 208938 64454 209494
rect 62288 187174 62608 187206
rect 62288 186938 62330 187174
rect 62566 186938 62608 187174
rect 62288 186854 62608 186938
rect 62288 186618 62330 186854
rect 62566 186618 62608 186854
rect 62288 186586 62608 186618
rect 60114 169218 60146 169774
rect 60702 169218 60734 169774
rect 60114 133774 60734 169218
rect 63834 173494 64454 208938
rect 63834 172938 63866 173494
rect 64422 172938 64454 173494
rect 62288 151174 62608 151206
rect 62288 150938 62330 151174
rect 62566 150938 62608 151174
rect 62288 150854 62608 150938
rect 62288 150618 62330 150854
rect 62566 150618 62608 150854
rect 62288 150586 62608 150618
rect 60114 133218 60146 133774
rect 60702 133218 60734 133774
rect 60114 97774 60734 133218
rect 63834 137494 64454 172938
rect 63834 136938 63866 137494
rect 64422 136938 64454 137494
rect 62288 115174 62608 115206
rect 62288 114938 62330 115174
rect 62566 114938 62608 115174
rect 62288 114854 62608 114938
rect 62288 114618 62330 114854
rect 62566 114618 62608 114854
rect 62288 114586 62608 114618
rect 60114 97218 60146 97774
rect 60702 97218 60734 97774
rect 60114 61774 60734 97218
rect 63834 101494 64454 136938
rect 63834 100938 63866 101494
rect 64422 100938 64454 101494
rect 62288 79174 62608 79206
rect 62288 78938 62330 79174
rect 62566 78938 62608 79174
rect 62288 78854 62608 78938
rect 62288 78618 62330 78854
rect 62566 78618 62608 78854
rect 62288 78586 62608 78618
rect 60114 61218 60146 61774
rect 60702 61218 60734 61774
rect 60114 25774 60734 61218
rect 63834 65494 64454 100938
rect 63834 64938 63866 65494
rect 64422 64938 64454 65494
rect 62288 43174 62608 43206
rect 62288 42938 62330 43174
rect 62566 42938 62608 43174
rect 62288 42854 62608 42938
rect 62288 42618 62330 42854
rect 62566 42618 62608 42854
rect 62288 42586 62608 42618
rect 60114 25218 60146 25774
rect 60702 25218 60734 25774
rect 59859 3908 59925 3909
rect 59859 3844 59860 3908
rect 59924 3844 59925 3908
rect 59859 3843 59925 3844
rect 59862 2821 59922 3843
rect 59859 2820 59925 2821
rect 59859 2756 59860 2820
rect 59924 2756 59925 2820
rect 59859 2755 59925 2756
rect 56394 -5702 56426 -5146
rect 56982 -5702 57014 -5146
rect 56394 -7654 57014 -5702
rect 60114 -6106 60734 25218
rect 63834 29494 64454 64938
rect 63834 28938 63866 29494
rect 64422 28938 64454 29494
rect 62288 7174 62608 7206
rect 62288 6938 62330 7174
rect 62566 6938 62608 7174
rect 62288 6854 62608 6938
rect 62288 6618 62330 6854
rect 62566 6618 62608 6854
rect 62288 6586 62608 6618
rect 60114 -6662 60146 -6106
rect 60702 -6662 60734 -6106
rect 60114 -7654 60734 -6662
rect 63834 -7066 64454 28938
rect 63834 -7622 63866 -7066
rect 64422 -7622 64454 -7066
rect 63834 -7654 64454 -7622
rect 73794 704838 74414 711590
rect 73794 704282 73826 704838
rect 74382 704282 74414 704838
rect 73794 687454 74414 704282
rect 73794 686898 73826 687454
rect 74382 686898 74414 687454
rect 73794 651454 74414 686898
rect 73794 650898 73826 651454
rect 74382 650898 74414 651454
rect 73794 615454 74414 650898
rect 73794 614898 73826 615454
rect 74382 614898 74414 615454
rect 73794 579454 74414 614898
rect 73794 578898 73826 579454
rect 74382 578898 74414 579454
rect 73794 543454 74414 578898
rect 73794 542898 73826 543454
rect 74382 542898 74414 543454
rect 73794 507454 74414 542898
rect 73794 506898 73826 507454
rect 74382 506898 74414 507454
rect 73794 471454 74414 506898
rect 73794 470898 73826 471454
rect 74382 470898 74414 471454
rect 73794 435454 74414 470898
rect 73794 434898 73826 435454
rect 74382 434898 74414 435454
rect 73794 399454 74414 434898
rect 73794 398898 73826 399454
rect 74382 398898 74414 399454
rect 73794 363454 74414 398898
rect 73794 362898 73826 363454
rect 74382 362898 74414 363454
rect 73794 327454 74414 362898
rect 77514 705798 78134 711590
rect 77514 705242 77546 705798
rect 78102 705242 78134 705798
rect 77514 691174 78134 705242
rect 77514 690618 77546 691174
rect 78102 690618 78134 691174
rect 77514 655174 78134 690618
rect 77514 654618 77546 655174
rect 78102 654618 78134 655174
rect 77514 619174 78134 654618
rect 77514 618618 77546 619174
rect 78102 618618 78134 619174
rect 77514 583174 78134 618618
rect 77514 582618 77546 583174
rect 78102 582618 78134 583174
rect 77514 547174 78134 582618
rect 77514 546618 77546 547174
rect 78102 546618 78134 547174
rect 77514 511174 78134 546618
rect 77514 510618 77546 511174
rect 78102 510618 78134 511174
rect 77514 475174 78134 510618
rect 77514 474618 77546 475174
rect 78102 474618 78134 475174
rect 77514 439174 78134 474618
rect 77514 438618 77546 439174
rect 78102 438618 78134 439174
rect 77514 403174 78134 438618
rect 77514 402618 77546 403174
rect 78102 402618 78134 403174
rect 77514 367174 78134 402618
rect 77514 366618 77546 367174
rect 78102 366618 78134 367174
rect 77514 354980 78134 366618
rect 81234 706758 81854 711590
rect 81234 706202 81266 706758
rect 81822 706202 81854 706758
rect 81234 694894 81854 706202
rect 81234 694338 81266 694894
rect 81822 694338 81854 694894
rect 81234 658894 81854 694338
rect 81234 658338 81266 658894
rect 81822 658338 81854 658894
rect 81234 622894 81854 658338
rect 81234 622338 81266 622894
rect 81822 622338 81854 622894
rect 81234 586894 81854 622338
rect 81234 586338 81266 586894
rect 81822 586338 81854 586894
rect 81234 550894 81854 586338
rect 81234 550338 81266 550894
rect 81822 550338 81854 550894
rect 81234 514894 81854 550338
rect 81234 514338 81266 514894
rect 81822 514338 81854 514894
rect 81234 478894 81854 514338
rect 81234 478338 81266 478894
rect 81822 478338 81854 478894
rect 81234 442894 81854 478338
rect 81234 442338 81266 442894
rect 81822 442338 81854 442894
rect 81234 406894 81854 442338
rect 81234 406338 81266 406894
rect 81822 406338 81854 406894
rect 81234 370894 81854 406338
rect 81234 370338 81266 370894
rect 81822 370338 81854 370894
rect 81234 334894 81854 370338
rect 81234 334338 81266 334894
rect 81822 334338 81854 334894
rect 73794 326898 73826 327454
rect 74382 326898 74414 327454
rect 73794 291454 74414 326898
rect 77648 327454 77968 327486
rect 77648 327218 77690 327454
rect 77926 327218 77968 327454
rect 77648 327134 77968 327218
rect 77648 326898 77690 327134
rect 77926 326898 77968 327134
rect 77648 326866 77968 326898
rect 81234 298894 81854 334338
rect 81234 298338 81266 298894
rect 81822 298338 81854 298894
rect 73794 290898 73826 291454
rect 74382 290898 74414 291454
rect 73794 255454 74414 290898
rect 77648 291454 77968 291486
rect 77648 291218 77690 291454
rect 77926 291218 77968 291454
rect 77648 291134 77968 291218
rect 77648 290898 77690 291134
rect 77926 290898 77968 291134
rect 77648 290866 77968 290898
rect 81234 262894 81854 298338
rect 81234 262338 81266 262894
rect 81822 262338 81854 262894
rect 73794 254898 73826 255454
rect 74382 254898 74414 255454
rect 73794 219454 74414 254898
rect 77648 255454 77968 255486
rect 77648 255218 77690 255454
rect 77926 255218 77968 255454
rect 77648 255134 77968 255218
rect 77648 254898 77690 255134
rect 77926 254898 77968 255134
rect 77648 254866 77968 254898
rect 81234 226894 81854 262338
rect 81234 226338 81266 226894
rect 81822 226338 81854 226894
rect 73794 218898 73826 219454
rect 74382 218898 74414 219454
rect 73794 183454 74414 218898
rect 77648 219454 77968 219486
rect 77648 219218 77690 219454
rect 77926 219218 77968 219454
rect 77648 219134 77968 219218
rect 77648 218898 77690 219134
rect 77926 218898 77968 219134
rect 77648 218866 77968 218898
rect 81234 190894 81854 226338
rect 81234 190338 81266 190894
rect 81822 190338 81854 190894
rect 73794 182898 73826 183454
rect 74382 182898 74414 183454
rect 73794 147454 74414 182898
rect 77648 183454 77968 183486
rect 77648 183218 77690 183454
rect 77926 183218 77968 183454
rect 77648 183134 77968 183218
rect 77648 182898 77690 183134
rect 77926 182898 77968 183134
rect 77648 182866 77968 182898
rect 81234 154894 81854 190338
rect 81234 154338 81266 154894
rect 81822 154338 81854 154894
rect 73794 146898 73826 147454
rect 74382 146898 74414 147454
rect 73794 111454 74414 146898
rect 77648 147454 77968 147486
rect 77648 147218 77690 147454
rect 77926 147218 77968 147454
rect 77648 147134 77968 147218
rect 77648 146898 77690 147134
rect 77926 146898 77968 147134
rect 77648 146866 77968 146898
rect 81234 118894 81854 154338
rect 81234 118338 81266 118894
rect 81822 118338 81854 118894
rect 73794 110898 73826 111454
rect 74382 110898 74414 111454
rect 73794 75454 74414 110898
rect 77648 111454 77968 111486
rect 77648 111218 77690 111454
rect 77926 111218 77968 111454
rect 77648 111134 77968 111218
rect 77648 110898 77690 111134
rect 77926 110898 77968 111134
rect 77648 110866 77968 110898
rect 81234 82894 81854 118338
rect 81234 82338 81266 82894
rect 81822 82338 81854 82894
rect 73794 74898 73826 75454
rect 74382 74898 74414 75454
rect 73794 39454 74414 74898
rect 77648 75454 77968 75486
rect 77648 75218 77690 75454
rect 77926 75218 77968 75454
rect 77648 75134 77968 75218
rect 77648 74898 77690 75134
rect 77926 74898 77968 75134
rect 77648 74866 77968 74898
rect 81234 46894 81854 82338
rect 81234 46338 81266 46894
rect 81822 46338 81854 46894
rect 73794 38898 73826 39454
rect 74382 38898 74414 39454
rect 73794 3454 74414 38898
rect 77648 39454 77968 39486
rect 77648 39218 77690 39454
rect 77926 39218 77968 39454
rect 77648 39134 77968 39218
rect 77648 38898 77690 39134
rect 77926 38898 77968 39134
rect 77648 38866 77968 38898
rect 73794 2898 73826 3454
rect 74382 2898 74414 3454
rect 73794 -346 74414 2898
rect 73794 -902 73826 -346
rect 74382 -902 74414 -346
rect 73794 -7654 74414 -902
rect 81234 10894 81854 46338
rect 81234 10338 81266 10894
rect 81822 10338 81854 10894
rect 81234 -2266 81854 10338
rect 81234 -2822 81266 -2266
rect 81822 -2822 81854 -2266
rect 81234 -7654 81854 -2822
rect 84954 707718 85574 711590
rect 84954 707162 84986 707718
rect 85542 707162 85574 707718
rect 84954 698614 85574 707162
rect 84954 698058 84986 698614
rect 85542 698058 85574 698614
rect 84954 662614 85574 698058
rect 84954 662058 84986 662614
rect 85542 662058 85574 662614
rect 84954 626614 85574 662058
rect 84954 626058 84986 626614
rect 85542 626058 85574 626614
rect 84954 590614 85574 626058
rect 84954 590058 84986 590614
rect 85542 590058 85574 590614
rect 84954 554614 85574 590058
rect 84954 554058 84986 554614
rect 85542 554058 85574 554614
rect 84954 518614 85574 554058
rect 84954 518058 84986 518614
rect 85542 518058 85574 518614
rect 84954 482614 85574 518058
rect 84954 482058 84986 482614
rect 85542 482058 85574 482614
rect 84954 446614 85574 482058
rect 84954 446058 84986 446614
rect 85542 446058 85574 446614
rect 84954 410614 85574 446058
rect 84954 410058 84986 410614
rect 85542 410058 85574 410614
rect 84954 374614 85574 410058
rect 84954 374058 84986 374614
rect 85542 374058 85574 374614
rect 84954 338614 85574 374058
rect 84954 338058 84986 338614
rect 85542 338058 85574 338614
rect 84954 302614 85574 338058
rect 84954 302058 84986 302614
rect 85542 302058 85574 302614
rect 84954 266614 85574 302058
rect 84954 266058 84986 266614
rect 85542 266058 85574 266614
rect 84954 230614 85574 266058
rect 84954 230058 84986 230614
rect 85542 230058 85574 230614
rect 84954 194614 85574 230058
rect 84954 194058 84986 194614
rect 85542 194058 85574 194614
rect 84954 158614 85574 194058
rect 84954 158058 84986 158614
rect 85542 158058 85574 158614
rect 84954 122614 85574 158058
rect 84954 122058 84986 122614
rect 85542 122058 85574 122614
rect 84954 86614 85574 122058
rect 84954 86058 84986 86614
rect 85542 86058 85574 86614
rect 84954 50614 85574 86058
rect 84954 50058 84986 50614
rect 85542 50058 85574 50614
rect 84954 14614 85574 50058
rect 84954 14058 84986 14614
rect 85542 14058 85574 14614
rect 84954 -3226 85574 14058
rect 84954 -3782 84986 -3226
rect 85542 -3782 85574 -3226
rect 84954 -7654 85574 -3782
rect 88674 708678 89294 711590
rect 88674 708122 88706 708678
rect 89262 708122 89294 708678
rect 88674 666334 89294 708122
rect 88674 665778 88706 666334
rect 89262 665778 89294 666334
rect 88674 630334 89294 665778
rect 88674 629778 88706 630334
rect 89262 629778 89294 630334
rect 88674 594334 89294 629778
rect 88674 593778 88706 594334
rect 89262 593778 89294 594334
rect 88674 558334 89294 593778
rect 88674 557778 88706 558334
rect 89262 557778 89294 558334
rect 88674 522334 89294 557778
rect 88674 521778 88706 522334
rect 89262 521778 89294 522334
rect 88674 486334 89294 521778
rect 88674 485778 88706 486334
rect 89262 485778 89294 486334
rect 88674 450334 89294 485778
rect 88674 449778 88706 450334
rect 89262 449778 89294 450334
rect 88674 414334 89294 449778
rect 88674 413778 88706 414334
rect 89262 413778 89294 414334
rect 88674 378334 89294 413778
rect 88674 377778 88706 378334
rect 89262 377778 89294 378334
rect 88674 342334 89294 377778
rect 92394 709638 93014 711590
rect 92394 709082 92426 709638
rect 92982 709082 93014 709638
rect 92394 670054 93014 709082
rect 92394 669498 92426 670054
rect 92982 669498 93014 670054
rect 92394 634054 93014 669498
rect 92394 633498 92426 634054
rect 92982 633498 93014 634054
rect 92394 598054 93014 633498
rect 92394 597498 92426 598054
rect 92982 597498 93014 598054
rect 92394 562054 93014 597498
rect 92394 561498 92426 562054
rect 92982 561498 93014 562054
rect 92394 526054 93014 561498
rect 92394 525498 92426 526054
rect 92982 525498 93014 526054
rect 92394 490054 93014 525498
rect 92394 489498 92426 490054
rect 92982 489498 93014 490054
rect 92394 454054 93014 489498
rect 92394 453498 92426 454054
rect 92982 453498 93014 454054
rect 92394 418054 93014 453498
rect 92394 417498 92426 418054
rect 92982 417498 93014 418054
rect 92394 382054 93014 417498
rect 92394 381498 92426 382054
rect 92982 381498 93014 382054
rect 92394 354980 93014 381498
rect 96114 710598 96734 711590
rect 96114 710042 96146 710598
rect 96702 710042 96734 710598
rect 96114 673774 96734 710042
rect 96114 673218 96146 673774
rect 96702 673218 96734 673774
rect 96114 637774 96734 673218
rect 96114 637218 96146 637774
rect 96702 637218 96734 637774
rect 96114 601774 96734 637218
rect 96114 601218 96146 601774
rect 96702 601218 96734 601774
rect 96114 565774 96734 601218
rect 96114 565218 96146 565774
rect 96702 565218 96734 565774
rect 96114 529774 96734 565218
rect 96114 529218 96146 529774
rect 96702 529218 96734 529774
rect 96114 493774 96734 529218
rect 96114 493218 96146 493774
rect 96702 493218 96734 493774
rect 96114 457774 96734 493218
rect 96114 457218 96146 457774
rect 96702 457218 96734 457774
rect 96114 421774 96734 457218
rect 96114 421218 96146 421774
rect 96702 421218 96734 421774
rect 96114 385774 96734 421218
rect 96114 385218 96146 385774
rect 96702 385218 96734 385774
rect 88674 341778 88706 342334
rect 89262 341778 89294 342334
rect 88674 306334 89294 341778
rect 96114 349774 96734 385218
rect 96114 349218 96146 349774
rect 96702 349218 96734 349774
rect 93008 331174 93328 331206
rect 93008 330938 93050 331174
rect 93286 330938 93328 331174
rect 93008 330854 93328 330938
rect 93008 330618 93050 330854
rect 93286 330618 93328 330854
rect 93008 330586 93328 330618
rect 88674 305778 88706 306334
rect 89262 305778 89294 306334
rect 88674 270334 89294 305778
rect 96114 313774 96734 349218
rect 96114 313218 96146 313774
rect 96702 313218 96734 313774
rect 93008 295174 93328 295206
rect 93008 294938 93050 295174
rect 93286 294938 93328 295174
rect 93008 294854 93328 294938
rect 93008 294618 93050 294854
rect 93286 294618 93328 294854
rect 93008 294586 93328 294618
rect 88674 269778 88706 270334
rect 89262 269778 89294 270334
rect 88674 234334 89294 269778
rect 96114 277774 96734 313218
rect 96114 277218 96146 277774
rect 96702 277218 96734 277774
rect 93008 259174 93328 259206
rect 93008 258938 93050 259174
rect 93286 258938 93328 259174
rect 93008 258854 93328 258938
rect 93008 258618 93050 258854
rect 93286 258618 93328 258854
rect 93008 258586 93328 258618
rect 88674 233778 88706 234334
rect 89262 233778 89294 234334
rect 88674 198334 89294 233778
rect 96114 241774 96734 277218
rect 96114 241218 96146 241774
rect 96702 241218 96734 241774
rect 93008 223174 93328 223206
rect 93008 222938 93050 223174
rect 93286 222938 93328 223174
rect 93008 222854 93328 222938
rect 93008 222618 93050 222854
rect 93286 222618 93328 222854
rect 93008 222586 93328 222618
rect 88674 197778 88706 198334
rect 89262 197778 89294 198334
rect 88674 162334 89294 197778
rect 96114 205774 96734 241218
rect 96114 205218 96146 205774
rect 96702 205218 96734 205774
rect 93008 187174 93328 187206
rect 93008 186938 93050 187174
rect 93286 186938 93328 187174
rect 93008 186854 93328 186938
rect 93008 186618 93050 186854
rect 93286 186618 93328 186854
rect 93008 186586 93328 186618
rect 88674 161778 88706 162334
rect 89262 161778 89294 162334
rect 88674 126334 89294 161778
rect 96114 169774 96734 205218
rect 96114 169218 96146 169774
rect 96702 169218 96734 169774
rect 93008 151174 93328 151206
rect 93008 150938 93050 151174
rect 93286 150938 93328 151174
rect 93008 150854 93328 150938
rect 93008 150618 93050 150854
rect 93286 150618 93328 150854
rect 93008 150586 93328 150618
rect 88674 125778 88706 126334
rect 89262 125778 89294 126334
rect 88674 90334 89294 125778
rect 96114 133774 96734 169218
rect 96114 133218 96146 133774
rect 96702 133218 96734 133774
rect 93008 115174 93328 115206
rect 93008 114938 93050 115174
rect 93286 114938 93328 115174
rect 93008 114854 93328 114938
rect 93008 114618 93050 114854
rect 93286 114618 93328 114854
rect 93008 114586 93328 114618
rect 88674 89778 88706 90334
rect 89262 89778 89294 90334
rect 88674 54334 89294 89778
rect 96114 97774 96734 133218
rect 96114 97218 96146 97774
rect 96702 97218 96734 97774
rect 93008 79174 93328 79206
rect 93008 78938 93050 79174
rect 93286 78938 93328 79174
rect 93008 78854 93328 78938
rect 93008 78618 93050 78854
rect 93286 78618 93328 78854
rect 93008 78586 93328 78618
rect 88674 53778 88706 54334
rect 89262 53778 89294 54334
rect 88674 18334 89294 53778
rect 96114 61774 96734 97218
rect 96114 61218 96146 61774
rect 96702 61218 96734 61774
rect 93008 43174 93328 43206
rect 93008 42938 93050 43174
rect 93286 42938 93328 43174
rect 93008 42854 93328 42938
rect 93008 42618 93050 42854
rect 93286 42618 93328 42854
rect 93008 42586 93328 42618
rect 88674 17778 88706 18334
rect 89262 17778 89294 18334
rect 88674 -4186 89294 17778
rect 96114 25774 96734 61218
rect 96114 25218 96146 25774
rect 96702 25218 96734 25774
rect 93008 7174 93328 7206
rect 93008 6938 93050 7174
rect 93286 6938 93328 7174
rect 93008 6854 93328 6938
rect 93008 6618 93050 6854
rect 93286 6618 93328 6854
rect 93008 6586 93328 6618
rect 88674 -4742 88706 -4186
rect 89262 -4742 89294 -4186
rect 88674 -7654 89294 -4742
rect 96114 -6106 96734 25218
rect 96114 -6662 96146 -6106
rect 96702 -6662 96734 -6106
rect 96114 -7654 96734 -6662
rect 99834 711558 100454 711590
rect 99834 711002 99866 711558
rect 100422 711002 100454 711558
rect 99834 677494 100454 711002
rect 99834 676938 99866 677494
rect 100422 676938 100454 677494
rect 99834 641494 100454 676938
rect 99834 640938 99866 641494
rect 100422 640938 100454 641494
rect 99834 605494 100454 640938
rect 99834 604938 99866 605494
rect 100422 604938 100454 605494
rect 99834 569494 100454 604938
rect 99834 568938 99866 569494
rect 100422 568938 100454 569494
rect 99834 533494 100454 568938
rect 99834 532938 99866 533494
rect 100422 532938 100454 533494
rect 99834 497494 100454 532938
rect 99834 496938 99866 497494
rect 100422 496938 100454 497494
rect 99834 461494 100454 496938
rect 99834 460938 99866 461494
rect 100422 460938 100454 461494
rect 99834 425494 100454 460938
rect 99834 424938 99866 425494
rect 100422 424938 100454 425494
rect 99834 389494 100454 424938
rect 99834 388938 99866 389494
rect 100422 388938 100454 389494
rect 99834 353494 100454 388938
rect 99834 352938 99866 353494
rect 100422 352938 100454 353494
rect 99834 317494 100454 352938
rect 109794 704838 110414 711590
rect 109794 704282 109826 704838
rect 110382 704282 110414 704838
rect 109794 687454 110414 704282
rect 109794 686898 109826 687454
rect 110382 686898 110414 687454
rect 109794 651454 110414 686898
rect 109794 650898 109826 651454
rect 110382 650898 110414 651454
rect 109794 615454 110414 650898
rect 109794 614898 109826 615454
rect 110382 614898 110414 615454
rect 109794 579454 110414 614898
rect 109794 578898 109826 579454
rect 110382 578898 110414 579454
rect 109794 543454 110414 578898
rect 109794 542898 109826 543454
rect 110382 542898 110414 543454
rect 109794 507454 110414 542898
rect 109794 506898 109826 507454
rect 110382 506898 110414 507454
rect 109794 471454 110414 506898
rect 109794 470898 109826 471454
rect 110382 470898 110414 471454
rect 109794 435454 110414 470898
rect 109794 434898 109826 435454
rect 110382 434898 110414 435454
rect 109794 399454 110414 434898
rect 109794 398898 109826 399454
rect 110382 398898 110414 399454
rect 109794 363454 110414 398898
rect 109794 362898 109826 363454
rect 110382 362898 110414 363454
rect 108368 327454 108688 327486
rect 108368 327218 108410 327454
rect 108646 327218 108688 327454
rect 108368 327134 108688 327218
rect 108368 326898 108410 327134
rect 108646 326898 108688 327134
rect 108368 326866 108688 326898
rect 109794 327454 110414 362898
rect 109794 326898 109826 327454
rect 110382 326898 110414 327454
rect 99834 316938 99866 317494
rect 100422 316938 100454 317494
rect 99834 281494 100454 316938
rect 108368 291454 108688 291486
rect 108368 291218 108410 291454
rect 108646 291218 108688 291454
rect 108368 291134 108688 291218
rect 108368 290898 108410 291134
rect 108646 290898 108688 291134
rect 108368 290866 108688 290898
rect 109794 291454 110414 326898
rect 109794 290898 109826 291454
rect 110382 290898 110414 291454
rect 99834 280938 99866 281494
rect 100422 280938 100454 281494
rect 99834 245494 100454 280938
rect 108368 255454 108688 255486
rect 108368 255218 108410 255454
rect 108646 255218 108688 255454
rect 108368 255134 108688 255218
rect 108368 254898 108410 255134
rect 108646 254898 108688 255134
rect 108368 254866 108688 254898
rect 109794 255454 110414 290898
rect 109794 254898 109826 255454
rect 110382 254898 110414 255454
rect 99834 244938 99866 245494
rect 100422 244938 100454 245494
rect 99834 209494 100454 244938
rect 108368 219454 108688 219486
rect 108368 219218 108410 219454
rect 108646 219218 108688 219454
rect 108368 219134 108688 219218
rect 108368 218898 108410 219134
rect 108646 218898 108688 219134
rect 108368 218866 108688 218898
rect 109794 219454 110414 254898
rect 109794 218898 109826 219454
rect 110382 218898 110414 219454
rect 99834 208938 99866 209494
rect 100422 208938 100454 209494
rect 99834 173494 100454 208938
rect 108368 183454 108688 183486
rect 108368 183218 108410 183454
rect 108646 183218 108688 183454
rect 108368 183134 108688 183218
rect 108368 182898 108410 183134
rect 108646 182898 108688 183134
rect 108368 182866 108688 182898
rect 109794 183454 110414 218898
rect 109794 182898 109826 183454
rect 110382 182898 110414 183454
rect 99834 172938 99866 173494
rect 100422 172938 100454 173494
rect 99834 137494 100454 172938
rect 108368 147454 108688 147486
rect 108368 147218 108410 147454
rect 108646 147218 108688 147454
rect 108368 147134 108688 147218
rect 108368 146898 108410 147134
rect 108646 146898 108688 147134
rect 108368 146866 108688 146898
rect 109794 147454 110414 182898
rect 109794 146898 109826 147454
rect 110382 146898 110414 147454
rect 99834 136938 99866 137494
rect 100422 136938 100454 137494
rect 99834 101494 100454 136938
rect 108368 111454 108688 111486
rect 108368 111218 108410 111454
rect 108646 111218 108688 111454
rect 108368 111134 108688 111218
rect 108368 110898 108410 111134
rect 108646 110898 108688 111134
rect 108368 110866 108688 110898
rect 109794 111454 110414 146898
rect 109794 110898 109826 111454
rect 110382 110898 110414 111454
rect 99834 100938 99866 101494
rect 100422 100938 100454 101494
rect 99834 65494 100454 100938
rect 108368 75454 108688 75486
rect 108368 75218 108410 75454
rect 108646 75218 108688 75454
rect 108368 75134 108688 75218
rect 108368 74898 108410 75134
rect 108646 74898 108688 75134
rect 108368 74866 108688 74898
rect 109794 75454 110414 110898
rect 109794 74898 109826 75454
rect 110382 74898 110414 75454
rect 99834 64938 99866 65494
rect 100422 64938 100454 65494
rect 99834 29494 100454 64938
rect 108368 39454 108688 39486
rect 108368 39218 108410 39454
rect 108646 39218 108688 39454
rect 108368 39134 108688 39218
rect 108368 38898 108410 39134
rect 108646 38898 108688 39134
rect 108368 38866 108688 38898
rect 109794 39454 110414 74898
rect 109794 38898 109826 39454
rect 110382 38898 110414 39454
rect 99834 28938 99866 29494
rect 100422 28938 100454 29494
rect 99834 -7066 100454 28938
rect 99834 -7622 99866 -7066
rect 100422 -7622 100454 -7066
rect 99834 -7654 100454 -7622
rect 109794 3454 110414 38898
rect 109794 2898 109826 3454
rect 110382 2898 110414 3454
rect 109794 -346 110414 2898
rect 109794 -902 109826 -346
rect 110382 -902 110414 -346
rect 109794 -7654 110414 -902
rect 113514 705798 114134 711590
rect 113514 705242 113546 705798
rect 114102 705242 114134 705798
rect 113514 691174 114134 705242
rect 113514 690618 113546 691174
rect 114102 690618 114134 691174
rect 113514 655174 114134 690618
rect 113514 654618 113546 655174
rect 114102 654618 114134 655174
rect 113514 619174 114134 654618
rect 113514 618618 113546 619174
rect 114102 618618 114134 619174
rect 113514 583174 114134 618618
rect 113514 582618 113546 583174
rect 114102 582618 114134 583174
rect 113514 547174 114134 582618
rect 113514 546618 113546 547174
rect 114102 546618 114134 547174
rect 113514 511174 114134 546618
rect 113514 510618 113546 511174
rect 114102 510618 114134 511174
rect 113514 475174 114134 510618
rect 113514 474618 113546 475174
rect 114102 474618 114134 475174
rect 113514 439174 114134 474618
rect 113514 438618 113546 439174
rect 114102 438618 114134 439174
rect 113514 403174 114134 438618
rect 113514 402618 113546 403174
rect 114102 402618 114134 403174
rect 113514 367174 114134 402618
rect 113514 366618 113546 367174
rect 114102 366618 114134 367174
rect 113514 331174 114134 366618
rect 113514 330618 113546 331174
rect 114102 330618 114134 331174
rect 113514 295174 114134 330618
rect 113514 294618 113546 295174
rect 114102 294618 114134 295174
rect 113514 259174 114134 294618
rect 113514 258618 113546 259174
rect 114102 258618 114134 259174
rect 113514 223174 114134 258618
rect 113514 222618 113546 223174
rect 114102 222618 114134 223174
rect 113514 187174 114134 222618
rect 113514 186618 113546 187174
rect 114102 186618 114134 187174
rect 113514 151174 114134 186618
rect 113514 150618 113546 151174
rect 114102 150618 114134 151174
rect 113514 115174 114134 150618
rect 113514 114618 113546 115174
rect 114102 114618 114134 115174
rect 113514 79174 114134 114618
rect 113514 78618 113546 79174
rect 114102 78618 114134 79174
rect 113514 43174 114134 78618
rect 113514 42618 113546 43174
rect 114102 42618 114134 43174
rect 113514 7174 114134 42618
rect 113514 6618 113546 7174
rect 114102 6618 114134 7174
rect 113514 -1306 114134 6618
rect 113514 -1862 113546 -1306
rect 114102 -1862 114134 -1306
rect 113514 -7654 114134 -1862
rect 117234 706758 117854 711590
rect 117234 706202 117266 706758
rect 117822 706202 117854 706758
rect 117234 694894 117854 706202
rect 117234 694338 117266 694894
rect 117822 694338 117854 694894
rect 117234 658894 117854 694338
rect 117234 658338 117266 658894
rect 117822 658338 117854 658894
rect 117234 622894 117854 658338
rect 117234 622338 117266 622894
rect 117822 622338 117854 622894
rect 117234 586894 117854 622338
rect 117234 586338 117266 586894
rect 117822 586338 117854 586894
rect 117234 550894 117854 586338
rect 117234 550338 117266 550894
rect 117822 550338 117854 550894
rect 117234 514894 117854 550338
rect 117234 514338 117266 514894
rect 117822 514338 117854 514894
rect 117234 478894 117854 514338
rect 117234 478338 117266 478894
rect 117822 478338 117854 478894
rect 117234 442894 117854 478338
rect 117234 442338 117266 442894
rect 117822 442338 117854 442894
rect 117234 406894 117854 442338
rect 117234 406338 117266 406894
rect 117822 406338 117854 406894
rect 117234 370894 117854 406338
rect 117234 370338 117266 370894
rect 117822 370338 117854 370894
rect 117234 334894 117854 370338
rect 117234 334338 117266 334894
rect 117822 334338 117854 334894
rect 117234 298894 117854 334338
rect 117234 298338 117266 298894
rect 117822 298338 117854 298894
rect 117234 262894 117854 298338
rect 117234 262338 117266 262894
rect 117822 262338 117854 262894
rect 117234 226894 117854 262338
rect 117234 226338 117266 226894
rect 117822 226338 117854 226894
rect 117234 190894 117854 226338
rect 117234 190338 117266 190894
rect 117822 190338 117854 190894
rect 117234 154894 117854 190338
rect 117234 154338 117266 154894
rect 117822 154338 117854 154894
rect 117234 118894 117854 154338
rect 117234 118338 117266 118894
rect 117822 118338 117854 118894
rect 117234 82894 117854 118338
rect 117234 82338 117266 82894
rect 117822 82338 117854 82894
rect 117234 46894 117854 82338
rect 117234 46338 117266 46894
rect 117822 46338 117854 46894
rect 117234 10894 117854 46338
rect 117234 10338 117266 10894
rect 117822 10338 117854 10894
rect 117234 -2266 117854 10338
rect 117234 -2822 117266 -2266
rect 117822 -2822 117854 -2266
rect 117234 -7654 117854 -2822
rect 120954 707718 121574 711590
rect 120954 707162 120986 707718
rect 121542 707162 121574 707718
rect 120954 698614 121574 707162
rect 120954 698058 120986 698614
rect 121542 698058 121574 698614
rect 120954 662614 121574 698058
rect 120954 662058 120986 662614
rect 121542 662058 121574 662614
rect 120954 626614 121574 662058
rect 120954 626058 120986 626614
rect 121542 626058 121574 626614
rect 120954 590614 121574 626058
rect 120954 590058 120986 590614
rect 121542 590058 121574 590614
rect 120954 554614 121574 590058
rect 120954 554058 120986 554614
rect 121542 554058 121574 554614
rect 120954 518614 121574 554058
rect 120954 518058 120986 518614
rect 121542 518058 121574 518614
rect 120954 482614 121574 518058
rect 120954 482058 120986 482614
rect 121542 482058 121574 482614
rect 120954 446614 121574 482058
rect 120954 446058 120986 446614
rect 121542 446058 121574 446614
rect 120954 410614 121574 446058
rect 120954 410058 120986 410614
rect 121542 410058 121574 410614
rect 120954 374614 121574 410058
rect 120954 374058 120986 374614
rect 121542 374058 121574 374614
rect 120954 338614 121574 374058
rect 120954 338058 120986 338614
rect 121542 338058 121574 338614
rect 120954 302614 121574 338058
rect 124674 708678 125294 711590
rect 124674 708122 124706 708678
rect 125262 708122 125294 708678
rect 124674 666334 125294 708122
rect 124674 665778 124706 666334
rect 125262 665778 125294 666334
rect 124674 630334 125294 665778
rect 124674 629778 124706 630334
rect 125262 629778 125294 630334
rect 124674 594334 125294 629778
rect 124674 593778 124706 594334
rect 125262 593778 125294 594334
rect 124674 558334 125294 593778
rect 124674 557778 124706 558334
rect 125262 557778 125294 558334
rect 124674 522334 125294 557778
rect 124674 521778 124706 522334
rect 125262 521778 125294 522334
rect 124674 486334 125294 521778
rect 124674 485778 124706 486334
rect 125262 485778 125294 486334
rect 124674 450334 125294 485778
rect 124674 449778 124706 450334
rect 125262 449778 125294 450334
rect 124674 414334 125294 449778
rect 124674 413778 124706 414334
rect 125262 413778 125294 414334
rect 124674 378334 125294 413778
rect 124674 377778 124706 378334
rect 125262 377778 125294 378334
rect 124674 342334 125294 377778
rect 124674 341778 124706 342334
rect 125262 341778 125294 342334
rect 123728 331174 124048 331206
rect 123728 330938 123770 331174
rect 124006 330938 124048 331174
rect 123728 330854 124048 330938
rect 123728 330618 123770 330854
rect 124006 330618 124048 330854
rect 123728 330586 124048 330618
rect 120954 302058 120986 302614
rect 121542 302058 121574 302614
rect 120954 266614 121574 302058
rect 124674 306334 125294 341778
rect 124674 305778 124706 306334
rect 125262 305778 125294 306334
rect 123728 295174 124048 295206
rect 123728 294938 123770 295174
rect 124006 294938 124048 295174
rect 123728 294854 124048 294938
rect 123728 294618 123770 294854
rect 124006 294618 124048 294854
rect 123728 294586 124048 294618
rect 120954 266058 120986 266614
rect 121542 266058 121574 266614
rect 120954 230614 121574 266058
rect 124674 270334 125294 305778
rect 124674 269778 124706 270334
rect 125262 269778 125294 270334
rect 123728 259174 124048 259206
rect 123728 258938 123770 259174
rect 124006 258938 124048 259174
rect 123728 258854 124048 258938
rect 123728 258618 123770 258854
rect 124006 258618 124048 258854
rect 123728 258586 124048 258618
rect 120954 230058 120986 230614
rect 121542 230058 121574 230614
rect 120954 194614 121574 230058
rect 124674 234334 125294 269778
rect 124674 233778 124706 234334
rect 125262 233778 125294 234334
rect 123728 223174 124048 223206
rect 123728 222938 123770 223174
rect 124006 222938 124048 223174
rect 123728 222854 124048 222938
rect 123728 222618 123770 222854
rect 124006 222618 124048 222854
rect 123728 222586 124048 222618
rect 120954 194058 120986 194614
rect 121542 194058 121574 194614
rect 120954 158614 121574 194058
rect 124674 198334 125294 233778
rect 124674 197778 124706 198334
rect 125262 197778 125294 198334
rect 123728 187174 124048 187206
rect 123728 186938 123770 187174
rect 124006 186938 124048 187174
rect 123728 186854 124048 186938
rect 123728 186618 123770 186854
rect 124006 186618 124048 186854
rect 123728 186586 124048 186618
rect 120954 158058 120986 158614
rect 121542 158058 121574 158614
rect 120954 122614 121574 158058
rect 124674 162334 125294 197778
rect 124674 161778 124706 162334
rect 125262 161778 125294 162334
rect 123728 151174 124048 151206
rect 123728 150938 123770 151174
rect 124006 150938 124048 151174
rect 123728 150854 124048 150938
rect 123728 150618 123770 150854
rect 124006 150618 124048 150854
rect 123728 150586 124048 150618
rect 120954 122058 120986 122614
rect 121542 122058 121574 122614
rect 120954 86614 121574 122058
rect 124674 126334 125294 161778
rect 124674 125778 124706 126334
rect 125262 125778 125294 126334
rect 123728 115174 124048 115206
rect 123728 114938 123770 115174
rect 124006 114938 124048 115174
rect 123728 114854 124048 114938
rect 123728 114618 123770 114854
rect 124006 114618 124048 114854
rect 123728 114586 124048 114618
rect 120954 86058 120986 86614
rect 121542 86058 121574 86614
rect 120954 50614 121574 86058
rect 124674 90334 125294 125778
rect 124674 89778 124706 90334
rect 125262 89778 125294 90334
rect 123728 79174 124048 79206
rect 123728 78938 123770 79174
rect 124006 78938 124048 79174
rect 123728 78854 124048 78938
rect 123728 78618 123770 78854
rect 124006 78618 124048 78854
rect 123728 78586 124048 78618
rect 120954 50058 120986 50614
rect 121542 50058 121574 50614
rect 120954 14614 121574 50058
rect 124674 54334 125294 89778
rect 124674 53778 124706 54334
rect 125262 53778 125294 54334
rect 123728 43174 124048 43206
rect 123728 42938 123770 43174
rect 124006 42938 124048 43174
rect 123728 42854 124048 42938
rect 123728 42618 123770 42854
rect 124006 42618 124048 42854
rect 123728 42586 124048 42618
rect 120954 14058 120986 14614
rect 121542 14058 121574 14614
rect 120954 -3226 121574 14058
rect 124674 18334 125294 53778
rect 124674 17778 124706 18334
rect 125262 17778 125294 18334
rect 123728 7174 124048 7206
rect 123728 6938 123770 7174
rect 124006 6938 124048 7174
rect 123728 6854 124048 6938
rect 123728 6618 123770 6854
rect 124006 6618 124048 6854
rect 123728 6586 124048 6618
rect 120954 -3782 120986 -3226
rect 121542 -3782 121574 -3226
rect 120954 -7654 121574 -3782
rect 124674 -4186 125294 17778
rect 124674 -4742 124706 -4186
rect 125262 -4742 125294 -4186
rect 124674 -7654 125294 -4742
rect 128394 709638 129014 711590
rect 128394 709082 128426 709638
rect 128982 709082 129014 709638
rect 128394 670054 129014 709082
rect 128394 669498 128426 670054
rect 128982 669498 129014 670054
rect 128394 634054 129014 669498
rect 128394 633498 128426 634054
rect 128982 633498 129014 634054
rect 128394 598054 129014 633498
rect 128394 597498 128426 598054
rect 128982 597498 129014 598054
rect 128394 562054 129014 597498
rect 128394 561498 128426 562054
rect 128982 561498 129014 562054
rect 128394 526054 129014 561498
rect 128394 525498 128426 526054
rect 128982 525498 129014 526054
rect 128394 490054 129014 525498
rect 128394 489498 128426 490054
rect 128982 489498 129014 490054
rect 128394 454054 129014 489498
rect 128394 453498 128426 454054
rect 128982 453498 129014 454054
rect 128394 418054 129014 453498
rect 128394 417498 128426 418054
rect 128982 417498 129014 418054
rect 128394 382054 129014 417498
rect 128394 381498 128426 382054
rect 128982 381498 129014 382054
rect 128394 346054 129014 381498
rect 128394 345498 128426 346054
rect 128982 345498 129014 346054
rect 128394 310054 129014 345498
rect 128394 309498 128426 310054
rect 128982 309498 129014 310054
rect 128394 274054 129014 309498
rect 128394 273498 128426 274054
rect 128982 273498 129014 274054
rect 128394 238054 129014 273498
rect 128394 237498 128426 238054
rect 128982 237498 129014 238054
rect 128394 202054 129014 237498
rect 128394 201498 128426 202054
rect 128982 201498 129014 202054
rect 128394 166054 129014 201498
rect 128394 165498 128426 166054
rect 128982 165498 129014 166054
rect 128394 130054 129014 165498
rect 128394 129498 128426 130054
rect 128982 129498 129014 130054
rect 128394 94054 129014 129498
rect 128394 93498 128426 94054
rect 128982 93498 129014 94054
rect 128394 58054 129014 93498
rect 128394 57498 128426 58054
rect 128982 57498 129014 58054
rect 128394 22054 129014 57498
rect 128394 21498 128426 22054
rect 128982 21498 129014 22054
rect 128394 -5146 129014 21498
rect 128394 -5702 128426 -5146
rect 128982 -5702 129014 -5146
rect 128394 -7654 129014 -5702
rect 132114 710598 132734 711590
rect 132114 710042 132146 710598
rect 132702 710042 132734 710598
rect 132114 673774 132734 710042
rect 132114 673218 132146 673774
rect 132702 673218 132734 673774
rect 132114 637774 132734 673218
rect 132114 637218 132146 637774
rect 132702 637218 132734 637774
rect 132114 601774 132734 637218
rect 132114 601218 132146 601774
rect 132702 601218 132734 601774
rect 132114 565774 132734 601218
rect 132114 565218 132146 565774
rect 132702 565218 132734 565774
rect 132114 529774 132734 565218
rect 132114 529218 132146 529774
rect 132702 529218 132734 529774
rect 132114 493774 132734 529218
rect 132114 493218 132146 493774
rect 132702 493218 132734 493774
rect 132114 457774 132734 493218
rect 132114 457218 132146 457774
rect 132702 457218 132734 457774
rect 132114 421774 132734 457218
rect 132114 421218 132146 421774
rect 132702 421218 132734 421774
rect 132114 385774 132734 421218
rect 132114 385218 132146 385774
rect 132702 385218 132734 385774
rect 132114 349774 132734 385218
rect 132114 349218 132146 349774
rect 132702 349218 132734 349774
rect 132114 313774 132734 349218
rect 132114 313218 132146 313774
rect 132702 313218 132734 313774
rect 132114 277774 132734 313218
rect 132114 277218 132146 277774
rect 132702 277218 132734 277774
rect 132114 241774 132734 277218
rect 132114 241218 132146 241774
rect 132702 241218 132734 241774
rect 132114 205774 132734 241218
rect 132114 205218 132146 205774
rect 132702 205218 132734 205774
rect 132114 169774 132734 205218
rect 132114 169218 132146 169774
rect 132702 169218 132734 169774
rect 132114 133774 132734 169218
rect 132114 133218 132146 133774
rect 132702 133218 132734 133774
rect 132114 97774 132734 133218
rect 132114 97218 132146 97774
rect 132702 97218 132734 97774
rect 132114 61774 132734 97218
rect 132114 61218 132146 61774
rect 132702 61218 132734 61774
rect 132114 25774 132734 61218
rect 132114 25218 132146 25774
rect 132702 25218 132734 25774
rect 132114 -6106 132734 25218
rect 132114 -6662 132146 -6106
rect 132702 -6662 132734 -6106
rect 132114 -7654 132734 -6662
rect 135834 711558 136454 711590
rect 135834 711002 135866 711558
rect 136422 711002 136454 711558
rect 135834 677494 136454 711002
rect 135834 676938 135866 677494
rect 136422 676938 136454 677494
rect 135834 641494 136454 676938
rect 135834 640938 135866 641494
rect 136422 640938 136454 641494
rect 135834 605494 136454 640938
rect 135834 604938 135866 605494
rect 136422 604938 136454 605494
rect 135834 569494 136454 604938
rect 135834 568938 135866 569494
rect 136422 568938 136454 569494
rect 135834 533494 136454 568938
rect 135834 532938 135866 533494
rect 136422 532938 136454 533494
rect 135834 497494 136454 532938
rect 135834 496938 135866 497494
rect 136422 496938 136454 497494
rect 135834 461494 136454 496938
rect 135834 460938 135866 461494
rect 136422 460938 136454 461494
rect 135834 425494 136454 460938
rect 135834 424938 135866 425494
rect 136422 424938 136454 425494
rect 135834 389494 136454 424938
rect 135834 388938 135866 389494
rect 136422 388938 136454 389494
rect 135834 353494 136454 388938
rect 135834 352938 135866 353494
rect 136422 352938 136454 353494
rect 135834 317494 136454 352938
rect 145794 704838 146414 711590
rect 145794 704282 145826 704838
rect 146382 704282 146414 704838
rect 145794 687454 146414 704282
rect 145794 686898 145826 687454
rect 146382 686898 146414 687454
rect 145794 651454 146414 686898
rect 145794 650898 145826 651454
rect 146382 650898 146414 651454
rect 145794 615454 146414 650898
rect 145794 614898 145826 615454
rect 146382 614898 146414 615454
rect 145794 579454 146414 614898
rect 145794 578898 145826 579454
rect 146382 578898 146414 579454
rect 145794 543454 146414 578898
rect 145794 542898 145826 543454
rect 146382 542898 146414 543454
rect 145794 507454 146414 542898
rect 145794 506898 145826 507454
rect 146382 506898 146414 507454
rect 145794 471454 146414 506898
rect 145794 470898 145826 471454
rect 146382 470898 146414 471454
rect 145794 435454 146414 470898
rect 145794 434898 145826 435454
rect 146382 434898 146414 435454
rect 145794 399454 146414 434898
rect 145794 398898 145826 399454
rect 146382 398898 146414 399454
rect 145794 363454 146414 398898
rect 145794 362898 145826 363454
rect 146382 362898 146414 363454
rect 139088 327454 139408 327486
rect 139088 327218 139130 327454
rect 139366 327218 139408 327454
rect 139088 327134 139408 327218
rect 139088 326898 139130 327134
rect 139366 326898 139408 327134
rect 139088 326866 139408 326898
rect 145794 327454 146414 362898
rect 145794 326898 145826 327454
rect 146382 326898 146414 327454
rect 135834 316938 135866 317494
rect 136422 316938 136454 317494
rect 135834 281494 136454 316938
rect 139088 291454 139408 291486
rect 139088 291218 139130 291454
rect 139366 291218 139408 291454
rect 139088 291134 139408 291218
rect 139088 290898 139130 291134
rect 139366 290898 139408 291134
rect 139088 290866 139408 290898
rect 145794 291454 146414 326898
rect 145794 290898 145826 291454
rect 146382 290898 146414 291454
rect 135834 280938 135866 281494
rect 136422 280938 136454 281494
rect 135834 245494 136454 280938
rect 139088 255454 139408 255486
rect 139088 255218 139130 255454
rect 139366 255218 139408 255454
rect 139088 255134 139408 255218
rect 139088 254898 139130 255134
rect 139366 254898 139408 255134
rect 139088 254866 139408 254898
rect 145794 255454 146414 290898
rect 145794 254898 145826 255454
rect 146382 254898 146414 255454
rect 135834 244938 135866 245494
rect 136422 244938 136454 245494
rect 135834 209494 136454 244938
rect 139088 219454 139408 219486
rect 139088 219218 139130 219454
rect 139366 219218 139408 219454
rect 139088 219134 139408 219218
rect 139088 218898 139130 219134
rect 139366 218898 139408 219134
rect 139088 218866 139408 218898
rect 145794 219454 146414 254898
rect 145794 218898 145826 219454
rect 146382 218898 146414 219454
rect 135834 208938 135866 209494
rect 136422 208938 136454 209494
rect 135834 173494 136454 208938
rect 139088 183454 139408 183486
rect 139088 183218 139130 183454
rect 139366 183218 139408 183454
rect 139088 183134 139408 183218
rect 139088 182898 139130 183134
rect 139366 182898 139408 183134
rect 139088 182866 139408 182898
rect 145794 183454 146414 218898
rect 145794 182898 145826 183454
rect 146382 182898 146414 183454
rect 135834 172938 135866 173494
rect 136422 172938 136454 173494
rect 135834 137494 136454 172938
rect 139088 147454 139408 147486
rect 139088 147218 139130 147454
rect 139366 147218 139408 147454
rect 139088 147134 139408 147218
rect 139088 146898 139130 147134
rect 139366 146898 139408 147134
rect 139088 146866 139408 146898
rect 145794 147454 146414 182898
rect 145794 146898 145826 147454
rect 146382 146898 146414 147454
rect 135834 136938 135866 137494
rect 136422 136938 136454 137494
rect 135834 101494 136454 136938
rect 139088 111454 139408 111486
rect 139088 111218 139130 111454
rect 139366 111218 139408 111454
rect 139088 111134 139408 111218
rect 139088 110898 139130 111134
rect 139366 110898 139408 111134
rect 139088 110866 139408 110898
rect 145794 111454 146414 146898
rect 145794 110898 145826 111454
rect 146382 110898 146414 111454
rect 135834 100938 135866 101494
rect 136422 100938 136454 101494
rect 135834 65494 136454 100938
rect 139088 75454 139408 75486
rect 139088 75218 139130 75454
rect 139366 75218 139408 75454
rect 139088 75134 139408 75218
rect 139088 74898 139130 75134
rect 139366 74898 139408 75134
rect 139088 74866 139408 74898
rect 145794 75454 146414 110898
rect 145794 74898 145826 75454
rect 146382 74898 146414 75454
rect 135834 64938 135866 65494
rect 136422 64938 136454 65494
rect 135834 29494 136454 64938
rect 139088 39454 139408 39486
rect 139088 39218 139130 39454
rect 139366 39218 139408 39454
rect 139088 39134 139408 39218
rect 139088 38898 139130 39134
rect 139366 38898 139408 39134
rect 139088 38866 139408 38898
rect 145794 39454 146414 74898
rect 145794 38898 145826 39454
rect 146382 38898 146414 39454
rect 135834 28938 135866 29494
rect 136422 28938 136454 29494
rect 135834 -7066 136454 28938
rect 135834 -7622 135866 -7066
rect 136422 -7622 136454 -7066
rect 135834 -7654 136454 -7622
rect 145794 3454 146414 38898
rect 145794 2898 145826 3454
rect 146382 2898 146414 3454
rect 145794 -346 146414 2898
rect 145794 -902 145826 -346
rect 146382 -902 146414 -346
rect 145794 -7654 146414 -902
rect 149514 705798 150134 711590
rect 149514 705242 149546 705798
rect 150102 705242 150134 705798
rect 149514 691174 150134 705242
rect 149514 690618 149546 691174
rect 150102 690618 150134 691174
rect 149514 655174 150134 690618
rect 149514 654618 149546 655174
rect 150102 654618 150134 655174
rect 149514 619174 150134 654618
rect 149514 618618 149546 619174
rect 150102 618618 150134 619174
rect 149514 583174 150134 618618
rect 149514 582618 149546 583174
rect 150102 582618 150134 583174
rect 149514 547174 150134 582618
rect 149514 546618 149546 547174
rect 150102 546618 150134 547174
rect 149514 511174 150134 546618
rect 149514 510618 149546 511174
rect 150102 510618 150134 511174
rect 149514 475174 150134 510618
rect 149514 474618 149546 475174
rect 150102 474618 150134 475174
rect 149514 439174 150134 474618
rect 149514 438618 149546 439174
rect 150102 438618 150134 439174
rect 149514 403174 150134 438618
rect 149514 402618 149546 403174
rect 150102 402618 150134 403174
rect 149514 367174 150134 402618
rect 149514 366618 149546 367174
rect 150102 366618 150134 367174
rect 149514 331174 150134 366618
rect 149514 330618 149546 331174
rect 150102 330618 150134 331174
rect 149514 295174 150134 330618
rect 149514 294618 149546 295174
rect 150102 294618 150134 295174
rect 149514 259174 150134 294618
rect 149514 258618 149546 259174
rect 150102 258618 150134 259174
rect 149514 223174 150134 258618
rect 149514 222618 149546 223174
rect 150102 222618 150134 223174
rect 149514 187174 150134 222618
rect 149514 186618 149546 187174
rect 150102 186618 150134 187174
rect 149514 151174 150134 186618
rect 149514 150618 149546 151174
rect 150102 150618 150134 151174
rect 149514 115174 150134 150618
rect 149514 114618 149546 115174
rect 150102 114618 150134 115174
rect 149514 79174 150134 114618
rect 149514 78618 149546 79174
rect 150102 78618 150134 79174
rect 149514 43174 150134 78618
rect 149514 42618 149546 43174
rect 150102 42618 150134 43174
rect 149514 7174 150134 42618
rect 149514 6618 149546 7174
rect 150102 6618 150134 7174
rect 149514 -1306 150134 6618
rect 149514 -1862 149546 -1306
rect 150102 -1862 150134 -1306
rect 149514 -7654 150134 -1862
rect 153234 706758 153854 711590
rect 153234 706202 153266 706758
rect 153822 706202 153854 706758
rect 153234 694894 153854 706202
rect 153234 694338 153266 694894
rect 153822 694338 153854 694894
rect 153234 658894 153854 694338
rect 153234 658338 153266 658894
rect 153822 658338 153854 658894
rect 153234 622894 153854 658338
rect 153234 622338 153266 622894
rect 153822 622338 153854 622894
rect 153234 586894 153854 622338
rect 153234 586338 153266 586894
rect 153822 586338 153854 586894
rect 153234 550894 153854 586338
rect 153234 550338 153266 550894
rect 153822 550338 153854 550894
rect 153234 514894 153854 550338
rect 153234 514338 153266 514894
rect 153822 514338 153854 514894
rect 153234 478894 153854 514338
rect 153234 478338 153266 478894
rect 153822 478338 153854 478894
rect 153234 442894 153854 478338
rect 153234 442338 153266 442894
rect 153822 442338 153854 442894
rect 153234 406894 153854 442338
rect 153234 406338 153266 406894
rect 153822 406338 153854 406894
rect 153234 370894 153854 406338
rect 153234 370338 153266 370894
rect 153822 370338 153854 370894
rect 153234 334894 153854 370338
rect 153234 334338 153266 334894
rect 153822 334338 153854 334894
rect 153234 298894 153854 334338
rect 156954 707718 157574 711590
rect 156954 707162 156986 707718
rect 157542 707162 157574 707718
rect 156954 698614 157574 707162
rect 156954 698058 156986 698614
rect 157542 698058 157574 698614
rect 156954 662614 157574 698058
rect 156954 662058 156986 662614
rect 157542 662058 157574 662614
rect 156954 626614 157574 662058
rect 156954 626058 156986 626614
rect 157542 626058 157574 626614
rect 156954 590614 157574 626058
rect 156954 590058 156986 590614
rect 157542 590058 157574 590614
rect 156954 554614 157574 590058
rect 156954 554058 156986 554614
rect 157542 554058 157574 554614
rect 156954 518614 157574 554058
rect 156954 518058 156986 518614
rect 157542 518058 157574 518614
rect 156954 482614 157574 518058
rect 156954 482058 156986 482614
rect 157542 482058 157574 482614
rect 156954 446614 157574 482058
rect 156954 446058 156986 446614
rect 157542 446058 157574 446614
rect 156954 410614 157574 446058
rect 156954 410058 156986 410614
rect 157542 410058 157574 410614
rect 156954 374614 157574 410058
rect 156954 374058 156986 374614
rect 157542 374058 157574 374614
rect 156954 338614 157574 374058
rect 156954 338058 156986 338614
rect 157542 338058 157574 338614
rect 154448 331174 154768 331206
rect 154448 330938 154490 331174
rect 154726 330938 154768 331174
rect 154448 330854 154768 330938
rect 154448 330618 154490 330854
rect 154726 330618 154768 330854
rect 154448 330586 154768 330618
rect 153234 298338 153266 298894
rect 153822 298338 153854 298894
rect 153234 262894 153854 298338
rect 156954 302614 157574 338058
rect 156954 302058 156986 302614
rect 157542 302058 157574 302614
rect 154448 295174 154768 295206
rect 154448 294938 154490 295174
rect 154726 294938 154768 295174
rect 154448 294854 154768 294938
rect 154448 294618 154490 294854
rect 154726 294618 154768 294854
rect 154448 294586 154768 294618
rect 153234 262338 153266 262894
rect 153822 262338 153854 262894
rect 153234 226894 153854 262338
rect 156954 266614 157574 302058
rect 156954 266058 156986 266614
rect 157542 266058 157574 266614
rect 154448 259174 154768 259206
rect 154448 258938 154490 259174
rect 154726 258938 154768 259174
rect 154448 258854 154768 258938
rect 154448 258618 154490 258854
rect 154726 258618 154768 258854
rect 154448 258586 154768 258618
rect 153234 226338 153266 226894
rect 153822 226338 153854 226894
rect 153234 190894 153854 226338
rect 156954 230614 157574 266058
rect 156954 230058 156986 230614
rect 157542 230058 157574 230614
rect 154448 223174 154768 223206
rect 154448 222938 154490 223174
rect 154726 222938 154768 223174
rect 154448 222854 154768 222938
rect 154448 222618 154490 222854
rect 154726 222618 154768 222854
rect 154448 222586 154768 222618
rect 153234 190338 153266 190894
rect 153822 190338 153854 190894
rect 153234 154894 153854 190338
rect 156954 194614 157574 230058
rect 156954 194058 156986 194614
rect 157542 194058 157574 194614
rect 154448 187174 154768 187206
rect 154448 186938 154490 187174
rect 154726 186938 154768 187174
rect 154448 186854 154768 186938
rect 154448 186618 154490 186854
rect 154726 186618 154768 186854
rect 154448 186586 154768 186618
rect 153234 154338 153266 154894
rect 153822 154338 153854 154894
rect 153234 118894 153854 154338
rect 156954 158614 157574 194058
rect 156954 158058 156986 158614
rect 157542 158058 157574 158614
rect 154448 151174 154768 151206
rect 154448 150938 154490 151174
rect 154726 150938 154768 151174
rect 154448 150854 154768 150938
rect 154448 150618 154490 150854
rect 154726 150618 154768 150854
rect 154448 150586 154768 150618
rect 153234 118338 153266 118894
rect 153822 118338 153854 118894
rect 153234 82894 153854 118338
rect 156954 122614 157574 158058
rect 156954 122058 156986 122614
rect 157542 122058 157574 122614
rect 154448 115174 154768 115206
rect 154448 114938 154490 115174
rect 154726 114938 154768 115174
rect 154448 114854 154768 114938
rect 154448 114618 154490 114854
rect 154726 114618 154768 114854
rect 154448 114586 154768 114618
rect 153234 82338 153266 82894
rect 153822 82338 153854 82894
rect 153234 46894 153854 82338
rect 156954 86614 157574 122058
rect 156954 86058 156986 86614
rect 157542 86058 157574 86614
rect 154448 79174 154768 79206
rect 154448 78938 154490 79174
rect 154726 78938 154768 79174
rect 154448 78854 154768 78938
rect 154448 78618 154490 78854
rect 154726 78618 154768 78854
rect 154448 78586 154768 78618
rect 153234 46338 153266 46894
rect 153822 46338 153854 46894
rect 153234 10894 153854 46338
rect 156954 50614 157574 86058
rect 156954 50058 156986 50614
rect 157542 50058 157574 50614
rect 154448 43174 154768 43206
rect 154448 42938 154490 43174
rect 154726 42938 154768 43174
rect 154448 42854 154768 42938
rect 154448 42618 154490 42854
rect 154726 42618 154768 42854
rect 154448 42586 154768 42618
rect 153234 10338 153266 10894
rect 153822 10338 153854 10894
rect 153234 -2266 153854 10338
rect 156954 14614 157574 50058
rect 156954 14058 156986 14614
rect 157542 14058 157574 14614
rect 154448 7174 154768 7206
rect 154448 6938 154490 7174
rect 154726 6938 154768 7174
rect 154448 6854 154768 6938
rect 154448 6618 154490 6854
rect 154726 6618 154768 6854
rect 154448 6586 154768 6618
rect 153234 -2822 153266 -2266
rect 153822 -2822 153854 -2266
rect 153234 -7654 153854 -2822
rect 156954 -3226 157574 14058
rect 156954 -3782 156986 -3226
rect 157542 -3782 157574 -3226
rect 156954 -7654 157574 -3782
rect 160674 708678 161294 711590
rect 160674 708122 160706 708678
rect 161262 708122 161294 708678
rect 160674 666334 161294 708122
rect 160674 665778 160706 666334
rect 161262 665778 161294 666334
rect 160674 630334 161294 665778
rect 160674 629778 160706 630334
rect 161262 629778 161294 630334
rect 160674 594334 161294 629778
rect 160674 593778 160706 594334
rect 161262 593778 161294 594334
rect 160674 558334 161294 593778
rect 160674 557778 160706 558334
rect 161262 557778 161294 558334
rect 160674 522334 161294 557778
rect 160674 521778 160706 522334
rect 161262 521778 161294 522334
rect 160674 486334 161294 521778
rect 160674 485778 160706 486334
rect 161262 485778 161294 486334
rect 160674 450334 161294 485778
rect 160674 449778 160706 450334
rect 161262 449778 161294 450334
rect 160674 414334 161294 449778
rect 160674 413778 160706 414334
rect 161262 413778 161294 414334
rect 160674 378334 161294 413778
rect 160674 377778 160706 378334
rect 161262 377778 161294 378334
rect 160674 342334 161294 377778
rect 160674 341778 160706 342334
rect 161262 341778 161294 342334
rect 160674 306334 161294 341778
rect 160674 305778 160706 306334
rect 161262 305778 161294 306334
rect 160674 270334 161294 305778
rect 160674 269778 160706 270334
rect 161262 269778 161294 270334
rect 160674 234334 161294 269778
rect 160674 233778 160706 234334
rect 161262 233778 161294 234334
rect 160674 198334 161294 233778
rect 160674 197778 160706 198334
rect 161262 197778 161294 198334
rect 160674 162334 161294 197778
rect 160674 161778 160706 162334
rect 161262 161778 161294 162334
rect 160674 126334 161294 161778
rect 160674 125778 160706 126334
rect 161262 125778 161294 126334
rect 160674 90334 161294 125778
rect 160674 89778 160706 90334
rect 161262 89778 161294 90334
rect 160674 54334 161294 89778
rect 160674 53778 160706 54334
rect 161262 53778 161294 54334
rect 160674 18334 161294 53778
rect 160674 17778 160706 18334
rect 161262 17778 161294 18334
rect 160674 -4186 161294 17778
rect 160674 -4742 160706 -4186
rect 161262 -4742 161294 -4186
rect 160674 -7654 161294 -4742
rect 164394 709638 165014 711590
rect 164394 709082 164426 709638
rect 164982 709082 165014 709638
rect 164394 670054 165014 709082
rect 164394 669498 164426 670054
rect 164982 669498 165014 670054
rect 164394 634054 165014 669498
rect 164394 633498 164426 634054
rect 164982 633498 165014 634054
rect 164394 598054 165014 633498
rect 164394 597498 164426 598054
rect 164982 597498 165014 598054
rect 164394 562054 165014 597498
rect 164394 561498 164426 562054
rect 164982 561498 165014 562054
rect 164394 526054 165014 561498
rect 164394 525498 164426 526054
rect 164982 525498 165014 526054
rect 164394 490054 165014 525498
rect 164394 489498 164426 490054
rect 164982 489498 165014 490054
rect 164394 454054 165014 489498
rect 164394 453498 164426 454054
rect 164982 453498 165014 454054
rect 164394 418054 165014 453498
rect 164394 417498 164426 418054
rect 164982 417498 165014 418054
rect 164394 382054 165014 417498
rect 164394 381498 164426 382054
rect 164982 381498 165014 382054
rect 164394 346054 165014 381498
rect 164394 345498 164426 346054
rect 164982 345498 165014 346054
rect 164394 310054 165014 345498
rect 164394 309498 164426 310054
rect 164982 309498 165014 310054
rect 164394 274054 165014 309498
rect 164394 273498 164426 274054
rect 164982 273498 165014 274054
rect 164394 238054 165014 273498
rect 164394 237498 164426 238054
rect 164982 237498 165014 238054
rect 164394 202054 165014 237498
rect 164394 201498 164426 202054
rect 164982 201498 165014 202054
rect 164394 166054 165014 201498
rect 164394 165498 164426 166054
rect 164982 165498 165014 166054
rect 164394 130054 165014 165498
rect 164394 129498 164426 130054
rect 164982 129498 165014 130054
rect 164394 94054 165014 129498
rect 164394 93498 164426 94054
rect 164982 93498 165014 94054
rect 164394 58054 165014 93498
rect 164394 57498 164426 58054
rect 164982 57498 165014 58054
rect 164394 22054 165014 57498
rect 164394 21498 164426 22054
rect 164982 21498 165014 22054
rect 164394 -5146 165014 21498
rect 164394 -5702 164426 -5146
rect 164982 -5702 165014 -5146
rect 164394 -7654 165014 -5702
rect 168114 710598 168734 711590
rect 168114 710042 168146 710598
rect 168702 710042 168734 710598
rect 168114 673774 168734 710042
rect 168114 673218 168146 673774
rect 168702 673218 168734 673774
rect 168114 637774 168734 673218
rect 168114 637218 168146 637774
rect 168702 637218 168734 637774
rect 168114 601774 168734 637218
rect 168114 601218 168146 601774
rect 168702 601218 168734 601774
rect 168114 565774 168734 601218
rect 168114 565218 168146 565774
rect 168702 565218 168734 565774
rect 168114 529774 168734 565218
rect 168114 529218 168146 529774
rect 168702 529218 168734 529774
rect 168114 493774 168734 529218
rect 168114 493218 168146 493774
rect 168702 493218 168734 493774
rect 168114 457774 168734 493218
rect 168114 457218 168146 457774
rect 168702 457218 168734 457774
rect 168114 421774 168734 457218
rect 168114 421218 168146 421774
rect 168702 421218 168734 421774
rect 168114 385774 168734 421218
rect 168114 385218 168146 385774
rect 168702 385218 168734 385774
rect 168114 349774 168734 385218
rect 168114 349218 168146 349774
rect 168702 349218 168734 349774
rect 168114 313774 168734 349218
rect 171834 711558 172454 711590
rect 171834 711002 171866 711558
rect 172422 711002 172454 711558
rect 171834 677494 172454 711002
rect 171834 676938 171866 677494
rect 172422 676938 172454 677494
rect 171834 641494 172454 676938
rect 171834 640938 171866 641494
rect 172422 640938 172454 641494
rect 171834 605494 172454 640938
rect 171834 604938 171866 605494
rect 172422 604938 172454 605494
rect 171834 569494 172454 604938
rect 171834 568938 171866 569494
rect 172422 568938 172454 569494
rect 171834 533494 172454 568938
rect 171834 532938 171866 533494
rect 172422 532938 172454 533494
rect 171834 497494 172454 532938
rect 171834 496938 171866 497494
rect 172422 496938 172454 497494
rect 171834 461494 172454 496938
rect 171834 460938 171866 461494
rect 172422 460938 172454 461494
rect 171834 425494 172454 460938
rect 171834 424938 171866 425494
rect 172422 424938 172454 425494
rect 171834 389494 172454 424938
rect 171834 388938 171866 389494
rect 172422 388938 172454 389494
rect 171834 353494 172454 388938
rect 171834 352938 171866 353494
rect 172422 352938 172454 353494
rect 169808 327454 170128 327486
rect 169808 327218 169850 327454
rect 170086 327218 170128 327454
rect 169808 327134 170128 327218
rect 169808 326898 169850 327134
rect 170086 326898 170128 327134
rect 169808 326866 170128 326898
rect 168114 313218 168146 313774
rect 168702 313218 168734 313774
rect 168114 277774 168734 313218
rect 171834 317494 172454 352938
rect 171834 316938 171866 317494
rect 172422 316938 172454 317494
rect 169808 291454 170128 291486
rect 169808 291218 169850 291454
rect 170086 291218 170128 291454
rect 169808 291134 170128 291218
rect 169808 290898 169850 291134
rect 170086 290898 170128 291134
rect 169808 290866 170128 290898
rect 168114 277218 168146 277774
rect 168702 277218 168734 277774
rect 168114 241774 168734 277218
rect 171834 281494 172454 316938
rect 171834 280938 171866 281494
rect 172422 280938 172454 281494
rect 169808 255454 170128 255486
rect 169808 255218 169850 255454
rect 170086 255218 170128 255454
rect 169808 255134 170128 255218
rect 169808 254898 169850 255134
rect 170086 254898 170128 255134
rect 169808 254866 170128 254898
rect 168114 241218 168146 241774
rect 168702 241218 168734 241774
rect 168114 205774 168734 241218
rect 171834 245494 172454 280938
rect 171834 244938 171866 245494
rect 172422 244938 172454 245494
rect 169808 219454 170128 219486
rect 169808 219218 169850 219454
rect 170086 219218 170128 219454
rect 169808 219134 170128 219218
rect 169808 218898 169850 219134
rect 170086 218898 170128 219134
rect 169808 218866 170128 218898
rect 168114 205218 168146 205774
rect 168702 205218 168734 205774
rect 168114 169774 168734 205218
rect 171834 209494 172454 244938
rect 171834 208938 171866 209494
rect 172422 208938 172454 209494
rect 169808 183454 170128 183486
rect 169808 183218 169850 183454
rect 170086 183218 170128 183454
rect 169808 183134 170128 183218
rect 169808 182898 169850 183134
rect 170086 182898 170128 183134
rect 169808 182866 170128 182898
rect 168114 169218 168146 169774
rect 168702 169218 168734 169774
rect 168114 133774 168734 169218
rect 171834 173494 172454 208938
rect 171834 172938 171866 173494
rect 172422 172938 172454 173494
rect 169808 147454 170128 147486
rect 169808 147218 169850 147454
rect 170086 147218 170128 147454
rect 169808 147134 170128 147218
rect 169808 146898 169850 147134
rect 170086 146898 170128 147134
rect 169808 146866 170128 146898
rect 168114 133218 168146 133774
rect 168702 133218 168734 133774
rect 168114 97774 168734 133218
rect 171834 137494 172454 172938
rect 171834 136938 171866 137494
rect 172422 136938 172454 137494
rect 169808 111454 170128 111486
rect 169808 111218 169850 111454
rect 170086 111218 170128 111454
rect 169808 111134 170128 111218
rect 169808 110898 169850 111134
rect 170086 110898 170128 111134
rect 169808 110866 170128 110898
rect 168114 97218 168146 97774
rect 168702 97218 168734 97774
rect 168114 61774 168734 97218
rect 171834 101494 172454 136938
rect 171834 100938 171866 101494
rect 172422 100938 172454 101494
rect 169808 75454 170128 75486
rect 169808 75218 169850 75454
rect 170086 75218 170128 75454
rect 169808 75134 170128 75218
rect 169808 74898 169850 75134
rect 170086 74898 170128 75134
rect 169808 74866 170128 74898
rect 168114 61218 168146 61774
rect 168702 61218 168734 61774
rect 168114 25774 168734 61218
rect 171834 65494 172454 100938
rect 171834 64938 171866 65494
rect 172422 64938 172454 65494
rect 169808 39454 170128 39486
rect 169808 39218 169850 39454
rect 170086 39218 170128 39454
rect 169808 39134 170128 39218
rect 169808 38898 169850 39134
rect 170086 38898 170128 39134
rect 169808 38866 170128 38898
rect 168114 25218 168146 25774
rect 168702 25218 168734 25774
rect 168114 -6106 168734 25218
rect 168114 -6662 168146 -6106
rect 168702 -6662 168734 -6106
rect 168114 -7654 168734 -6662
rect 171834 29494 172454 64938
rect 171834 28938 171866 29494
rect 172422 28938 172454 29494
rect 171834 -7066 172454 28938
rect 171834 -7622 171866 -7066
rect 172422 -7622 172454 -7066
rect 171834 -7654 172454 -7622
rect 181794 704838 182414 711590
rect 181794 704282 181826 704838
rect 182382 704282 182414 704838
rect 181794 687454 182414 704282
rect 181794 686898 181826 687454
rect 182382 686898 182414 687454
rect 181794 651454 182414 686898
rect 181794 650898 181826 651454
rect 182382 650898 182414 651454
rect 181794 615454 182414 650898
rect 181794 614898 181826 615454
rect 182382 614898 182414 615454
rect 181794 579454 182414 614898
rect 181794 578898 181826 579454
rect 182382 578898 182414 579454
rect 181794 543454 182414 578898
rect 181794 542898 181826 543454
rect 182382 542898 182414 543454
rect 181794 507454 182414 542898
rect 181794 506898 181826 507454
rect 182382 506898 182414 507454
rect 181794 471454 182414 506898
rect 181794 470898 181826 471454
rect 182382 470898 182414 471454
rect 181794 435454 182414 470898
rect 181794 434898 181826 435454
rect 182382 434898 182414 435454
rect 181794 399454 182414 434898
rect 181794 398898 181826 399454
rect 182382 398898 182414 399454
rect 181794 363454 182414 398898
rect 181794 362898 181826 363454
rect 182382 362898 182414 363454
rect 181794 327454 182414 362898
rect 185514 705798 186134 711590
rect 185514 705242 185546 705798
rect 186102 705242 186134 705798
rect 185514 691174 186134 705242
rect 185514 690618 185546 691174
rect 186102 690618 186134 691174
rect 185514 655174 186134 690618
rect 185514 654618 185546 655174
rect 186102 654618 186134 655174
rect 185514 619174 186134 654618
rect 185514 618618 185546 619174
rect 186102 618618 186134 619174
rect 185514 583174 186134 618618
rect 185514 582618 185546 583174
rect 186102 582618 186134 583174
rect 185514 547174 186134 582618
rect 185514 546618 185546 547174
rect 186102 546618 186134 547174
rect 185514 511174 186134 546618
rect 185514 510618 185546 511174
rect 186102 510618 186134 511174
rect 185514 475174 186134 510618
rect 185514 474618 185546 475174
rect 186102 474618 186134 475174
rect 185514 439174 186134 474618
rect 185514 438618 185546 439174
rect 186102 438618 186134 439174
rect 185514 403174 186134 438618
rect 185514 402618 185546 403174
rect 186102 402618 186134 403174
rect 185514 367174 186134 402618
rect 185514 366618 185546 367174
rect 186102 366618 186134 367174
rect 185514 354980 186134 366618
rect 189234 706758 189854 711590
rect 189234 706202 189266 706758
rect 189822 706202 189854 706758
rect 189234 694894 189854 706202
rect 189234 694338 189266 694894
rect 189822 694338 189854 694894
rect 189234 658894 189854 694338
rect 189234 658338 189266 658894
rect 189822 658338 189854 658894
rect 189234 622894 189854 658338
rect 189234 622338 189266 622894
rect 189822 622338 189854 622894
rect 189234 586894 189854 622338
rect 189234 586338 189266 586894
rect 189822 586338 189854 586894
rect 189234 550894 189854 586338
rect 189234 550338 189266 550894
rect 189822 550338 189854 550894
rect 189234 514894 189854 550338
rect 189234 514338 189266 514894
rect 189822 514338 189854 514894
rect 189234 478894 189854 514338
rect 189234 478338 189266 478894
rect 189822 478338 189854 478894
rect 189234 442894 189854 478338
rect 189234 442338 189266 442894
rect 189822 442338 189854 442894
rect 189234 406894 189854 442338
rect 189234 406338 189266 406894
rect 189822 406338 189854 406894
rect 189234 370894 189854 406338
rect 189234 370338 189266 370894
rect 189822 370338 189854 370894
rect 189234 334894 189854 370338
rect 189234 334338 189266 334894
rect 189822 334338 189854 334894
rect 185168 331174 185488 331206
rect 185168 330938 185210 331174
rect 185446 330938 185488 331174
rect 185168 330854 185488 330938
rect 185168 330618 185210 330854
rect 185446 330618 185488 330854
rect 185168 330586 185488 330618
rect 181794 326898 181826 327454
rect 182382 326898 182414 327454
rect 181794 291454 182414 326898
rect 189234 298894 189854 334338
rect 189234 298338 189266 298894
rect 189822 298338 189854 298894
rect 185168 295174 185488 295206
rect 185168 294938 185210 295174
rect 185446 294938 185488 295174
rect 185168 294854 185488 294938
rect 185168 294618 185210 294854
rect 185446 294618 185488 294854
rect 185168 294586 185488 294618
rect 181794 290898 181826 291454
rect 182382 290898 182414 291454
rect 181794 255454 182414 290898
rect 189234 262894 189854 298338
rect 189234 262338 189266 262894
rect 189822 262338 189854 262894
rect 185168 259174 185488 259206
rect 185168 258938 185210 259174
rect 185446 258938 185488 259174
rect 185168 258854 185488 258938
rect 185168 258618 185210 258854
rect 185446 258618 185488 258854
rect 185168 258586 185488 258618
rect 181794 254898 181826 255454
rect 182382 254898 182414 255454
rect 181794 219454 182414 254898
rect 189234 226894 189854 262338
rect 189234 226338 189266 226894
rect 189822 226338 189854 226894
rect 185168 223174 185488 223206
rect 185168 222938 185210 223174
rect 185446 222938 185488 223174
rect 185168 222854 185488 222938
rect 185168 222618 185210 222854
rect 185446 222618 185488 222854
rect 185168 222586 185488 222618
rect 181794 218898 181826 219454
rect 182382 218898 182414 219454
rect 181794 183454 182414 218898
rect 189234 190894 189854 226338
rect 189234 190338 189266 190894
rect 189822 190338 189854 190894
rect 185168 187174 185488 187206
rect 185168 186938 185210 187174
rect 185446 186938 185488 187174
rect 185168 186854 185488 186938
rect 185168 186618 185210 186854
rect 185446 186618 185488 186854
rect 185168 186586 185488 186618
rect 181794 182898 181826 183454
rect 182382 182898 182414 183454
rect 181794 147454 182414 182898
rect 189234 154894 189854 190338
rect 189234 154338 189266 154894
rect 189822 154338 189854 154894
rect 185168 151174 185488 151206
rect 185168 150938 185210 151174
rect 185446 150938 185488 151174
rect 185168 150854 185488 150938
rect 185168 150618 185210 150854
rect 185446 150618 185488 150854
rect 185168 150586 185488 150618
rect 181794 146898 181826 147454
rect 182382 146898 182414 147454
rect 181794 111454 182414 146898
rect 189234 118894 189854 154338
rect 189234 118338 189266 118894
rect 189822 118338 189854 118894
rect 185168 115174 185488 115206
rect 185168 114938 185210 115174
rect 185446 114938 185488 115174
rect 185168 114854 185488 114938
rect 185168 114618 185210 114854
rect 185446 114618 185488 114854
rect 185168 114586 185488 114618
rect 181794 110898 181826 111454
rect 182382 110898 182414 111454
rect 181794 75454 182414 110898
rect 189234 82894 189854 118338
rect 189234 82338 189266 82894
rect 189822 82338 189854 82894
rect 185168 79174 185488 79206
rect 185168 78938 185210 79174
rect 185446 78938 185488 79174
rect 185168 78854 185488 78938
rect 185168 78618 185210 78854
rect 185446 78618 185488 78854
rect 185168 78586 185488 78618
rect 181794 74898 181826 75454
rect 182382 74898 182414 75454
rect 181794 39454 182414 74898
rect 189234 46894 189854 82338
rect 189234 46338 189266 46894
rect 189822 46338 189854 46894
rect 185168 43174 185488 43206
rect 185168 42938 185210 43174
rect 185446 42938 185488 43174
rect 185168 42854 185488 42938
rect 185168 42618 185210 42854
rect 185446 42618 185488 42854
rect 185168 42586 185488 42618
rect 181794 38898 181826 39454
rect 182382 38898 182414 39454
rect 181794 3454 182414 38898
rect 189234 10894 189854 46338
rect 189234 10338 189266 10894
rect 189822 10338 189854 10894
rect 185168 7174 185488 7206
rect 185168 6938 185210 7174
rect 185446 6938 185488 7174
rect 185168 6854 185488 6938
rect 185168 6618 185210 6854
rect 185446 6618 185488 6854
rect 185168 6586 185488 6618
rect 181794 2898 181826 3454
rect 182382 2898 182414 3454
rect 181794 -346 182414 2898
rect 181794 -902 181826 -346
rect 182382 -902 182414 -346
rect 181794 -7654 182414 -902
rect 189234 -2266 189854 10338
rect 189234 -2822 189266 -2266
rect 189822 -2822 189854 -2266
rect 189234 -7654 189854 -2822
rect 192954 707718 193574 711590
rect 192954 707162 192986 707718
rect 193542 707162 193574 707718
rect 192954 698614 193574 707162
rect 192954 698058 192986 698614
rect 193542 698058 193574 698614
rect 192954 662614 193574 698058
rect 192954 662058 192986 662614
rect 193542 662058 193574 662614
rect 192954 626614 193574 662058
rect 192954 626058 192986 626614
rect 193542 626058 193574 626614
rect 192954 590614 193574 626058
rect 192954 590058 192986 590614
rect 193542 590058 193574 590614
rect 192954 554614 193574 590058
rect 192954 554058 192986 554614
rect 193542 554058 193574 554614
rect 192954 518614 193574 554058
rect 192954 518058 192986 518614
rect 193542 518058 193574 518614
rect 192954 482614 193574 518058
rect 192954 482058 192986 482614
rect 193542 482058 193574 482614
rect 192954 446614 193574 482058
rect 192954 446058 192986 446614
rect 193542 446058 193574 446614
rect 192954 410614 193574 446058
rect 192954 410058 192986 410614
rect 193542 410058 193574 410614
rect 192954 374614 193574 410058
rect 192954 374058 192986 374614
rect 193542 374058 193574 374614
rect 192954 338614 193574 374058
rect 192954 338058 192986 338614
rect 193542 338058 193574 338614
rect 192954 302614 193574 338058
rect 192954 302058 192986 302614
rect 193542 302058 193574 302614
rect 192954 266614 193574 302058
rect 192954 266058 192986 266614
rect 193542 266058 193574 266614
rect 192954 230614 193574 266058
rect 192954 230058 192986 230614
rect 193542 230058 193574 230614
rect 192954 194614 193574 230058
rect 192954 194058 192986 194614
rect 193542 194058 193574 194614
rect 192954 158614 193574 194058
rect 192954 158058 192986 158614
rect 193542 158058 193574 158614
rect 192954 122614 193574 158058
rect 192954 122058 192986 122614
rect 193542 122058 193574 122614
rect 192954 86614 193574 122058
rect 192954 86058 192986 86614
rect 193542 86058 193574 86614
rect 192954 50614 193574 86058
rect 192954 50058 192986 50614
rect 193542 50058 193574 50614
rect 192954 14614 193574 50058
rect 192954 14058 192986 14614
rect 193542 14058 193574 14614
rect 192954 -3226 193574 14058
rect 192954 -3782 192986 -3226
rect 193542 -3782 193574 -3226
rect 192954 -7654 193574 -3782
rect 196674 708678 197294 711590
rect 196674 708122 196706 708678
rect 197262 708122 197294 708678
rect 196674 666334 197294 708122
rect 196674 665778 196706 666334
rect 197262 665778 197294 666334
rect 196674 630334 197294 665778
rect 196674 629778 196706 630334
rect 197262 629778 197294 630334
rect 196674 594334 197294 629778
rect 196674 593778 196706 594334
rect 197262 593778 197294 594334
rect 196674 558334 197294 593778
rect 196674 557778 196706 558334
rect 197262 557778 197294 558334
rect 196674 522334 197294 557778
rect 196674 521778 196706 522334
rect 197262 521778 197294 522334
rect 196674 486334 197294 521778
rect 196674 485778 196706 486334
rect 197262 485778 197294 486334
rect 196674 450334 197294 485778
rect 196674 449778 196706 450334
rect 197262 449778 197294 450334
rect 196674 414334 197294 449778
rect 196674 413778 196706 414334
rect 197262 413778 197294 414334
rect 196674 378334 197294 413778
rect 196674 377778 196706 378334
rect 197262 377778 197294 378334
rect 196674 342334 197294 377778
rect 200394 709638 201014 711590
rect 200394 709082 200426 709638
rect 200982 709082 201014 709638
rect 200394 670054 201014 709082
rect 200394 669498 200426 670054
rect 200982 669498 201014 670054
rect 200394 634054 201014 669498
rect 200394 633498 200426 634054
rect 200982 633498 201014 634054
rect 200394 598054 201014 633498
rect 200394 597498 200426 598054
rect 200982 597498 201014 598054
rect 200394 562054 201014 597498
rect 200394 561498 200426 562054
rect 200982 561498 201014 562054
rect 200394 526054 201014 561498
rect 200394 525498 200426 526054
rect 200982 525498 201014 526054
rect 200394 490054 201014 525498
rect 200394 489498 200426 490054
rect 200982 489498 201014 490054
rect 200394 454054 201014 489498
rect 200394 453498 200426 454054
rect 200982 453498 201014 454054
rect 200394 418054 201014 453498
rect 200394 417498 200426 418054
rect 200982 417498 201014 418054
rect 200394 382054 201014 417498
rect 200394 381498 200426 382054
rect 200982 381498 201014 382054
rect 200394 354980 201014 381498
rect 204114 710598 204734 711590
rect 204114 710042 204146 710598
rect 204702 710042 204734 710598
rect 204114 673774 204734 710042
rect 204114 673218 204146 673774
rect 204702 673218 204734 673774
rect 204114 637774 204734 673218
rect 204114 637218 204146 637774
rect 204702 637218 204734 637774
rect 204114 601774 204734 637218
rect 204114 601218 204146 601774
rect 204702 601218 204734 601774
rect 204114 565774 204734 601218
rect 204114 565218 204146 565774
rect 204702 565218 204734 565774
rect 204114 529774 204734 565218
rect 204114 529218 204146 529774
rect 204702 529218 204734 529774
rect 204114 493774 204734 529218
rect 204114 493218 204146 493774
rect 204702 493218 204734 493774
rect 204114 457774 204734 493218
rect 204114 457218 204146 457774
rect 204702 457218 204734 457774
rect 204114 421774 204734 457218
rect 204114 421218 204146 421774
rect 204702 421218 204734 421774
rect 204114 385774 204734 421218
rect 204114 385218 204146 385774
rect 204702 385218 204734 385774
rect 196674 341778 196706 342334
rect 197262 341778 197294 342334
rect 196674 306334 197294 341778
rect 204114 349774 204734 385218
rect 204114 349218 204146 349774
rect 204702 349218 204734 349774
rect 200528 327454 200848 327486
rect 200528 327218 200570 327454
rect 200806 327218 200848 327454
rect 200528 327134 200848 327218
rect 200528 326898 200570 327134
rect 200806 326898 200848 327134
rect 200528 326866 200848 326898
rect 196674 305778 196706 306334
rect 197262 305778 197294 306334
rect 196674 270334 197294 305778
rect 204114 313774 204734 349218
rect 204114 313218 204146 313774
rect 204702 313218 204734 313774
rect 200528 291454 200848 291486
rect 200528 291218 200570 291454
rect 200806 291218 200848 291454
rect 200528 291134 200848 291218
rect 200528 290898 200570 291134
rect 200806 290898 200848 291134
rect 200528 290866 200848 290898
rect 196674 269778 196706 270334
rect 197262 269778 197294 270334
rect 196674 234334 197294 269778
rect 204114 277774 204734 313218
rect 204114 277218 204146 277774
rect 204702 277218 204734 277774
rect 200528 255454 200848 255486
rect 200528 255218 200570 255454
rect 200806 255218 200848 255454
rect 200528 255134 200848 255218
rect 200528 254898 200570 255134
rect 200806 254898 200848 255134
rect 200528 254866 200848 254898
rect 196674 233778 196706 234334
rect 197262 233778 197294 234334
rect 196674 198334 197294 233778
rect 204114 241774 204734 277218
rect 204114 241218 204146 241774
rect 204702 241218 204734 241774
rect 200528 219454 200848 219486
rect 200528 219218 200570 219454
rect 200806 219218 200848 219454
rect 200528 219134 200848 219218
rect 200528 218898 200570 219134
rect 200806 218898 200848 219134
rect 200528 218866 200848 218898
rect 196674 197778 196706 198334
rect 197262 197778 197294 198334
rect 196674 162334 197294 197778
rect 204114 205774 204734 241218
rect 204114 205218 204146 205774
rect 204702 205218 204734 205774
rect 200528 183454 200848 183486
rect 200528 183218 200570 183454
rect 200806 183218 200848 183454
rect 200528 183134 200848 183218
rect 200528 182898 200570 183134
rect 200806 182898 200848 183134
rect 200528 182866 200848 182898
rect 196674 161778 196706 162334
rect 197262 161778 197294 162334
rect 196674 126334 197294 161778
rect 204114 169774 204734 205218
rect 204114 169218 204146 169774
rect 204702 169218 204734 169774
rect 200528 147454 200848 147486
rect 200528 147218 200570 147454
rect 200806 147218 200848 147454
rect 200528 147134 200848 147218
rect 200528 146898 200570 147134
rect 200806 146898 200848 147134
rect 200528 146866 200848 146898
rect 196674 125778 196706 126334
rect 197262 125778 197294 126334
rect 196674 90334 197294 125778
rect 204114 133774 204734 169218
rect 204114 133218 204146 133774
rect 204702 133218 204734 133774
rect 200528 111454 200848 111486
rect 200528 111218 200570 111454
rect 200806 111218 200848 111454
rect 200528 111134 200848 111218
rect 200528 110898 200570 111134
rect 200806 110898 200848 111134
rect 200528 110866 200848 110898
rect 196674 89778 196706 90334
rect 197262 89778 197294 90334
rect 196674 54334 197294 89778
rect 204114 97774 204734 133218
rect 204114 97218 204146 97774
rect 204702 97218 204734 97774
rect 200528 75454 200848 75486
rect 200528 75218 200570 75454
rect 200806 75218 200848 75454
rect 200528 75134 200848 75218
rect 200528 74898 200570 75134
rect 200806 74898 200848 75134
rect 200528 74866 200848 74898
rect 196674 53778 196706 54334
rect 197262 53778 197294 54334
rect 196674 18334 197294 53778
rect 204114 61774 204734 97218
rect 204114 61218 204146 61774
rect 204702 61218 204734 61774
rect 200528 39454 200848 39486
rect 200528 39218 200570 39454
rect 200806 39218 200848 39454
rect 200528 39134 200848 39218
rect 200528 38898 200570 39134
rect 200806 38898 200848 39134
rect 200528 38866 200848 38898
rect 196674 17778 196706 18334
rect 197262 17778 197294 18334
rect 196674 -4186 197294 17778
rect 196674 -4742 196706 -4186
rect 197262 -4742 197294 -4186
rect 196674 -7654 197294 -4742
rect 204114 25774 204734 61218
rect 204114 25218 204146 25774
rect 204702 25218 204734 25774
rect 204114 -6106 204734 25218
rect 204114 -6662 204146 -6106
rect 204702 -6662 204734 -6106
rect 204114 -7654 204734 -6662
rect 207834 711558 208454 711590
rect 207834 711002 207866 711558
rect 208422 711002 208454 711558
rect 207834 677494 208454 711002
rect 207834 676938 207866 677494
rect 208422 676938 208454 677494
rect 207834 641494 208454 676938
rect 207834 640938 207866 641494
rect 208422 640938 208454 641494
rect 207834 605494 208454 640938
rect 207834 604938 207866 605494
rect 208422 604938 208454 605494
rect 207834 569494 208454 604938
rect 207834 568938 207866 569494
rect 208422 568938 208454 569494
rect 207834 533494 208454 568938
rect 207834 532938 207866 533494
rect 208422 532938 208454 533494
rect 207834 497494 208454 532938
rect 207834 496938 207866 497494
rect 208422 496938 208454 497494
rect 207834 461494 208454 496938
rect 207834 460938 207866 461494
rect 208422 460938 208454 461494
rect 207834 425494 208454 460938
rect 207834 424938 207866 425494
rect 208422 424938 208454 425494
rect 207834 389494 208454 424938
rect 207834 388938 207866 389494
rect 208422 388938 208454 389494
rect 207834 353494 208454 388938
rect 207834 352938 207866 353494
rect 208422 352938 208454 353494
rect 207834 317494 208454 352938
rect 217794 704838 218414 711590
rect 217794 704282 217826 704838
rect 218382 704282 218414 704838
rect 217794 687454 218414 704282
rect 217794 686898 217826 687454
rect 218382 686898 218414 687454
rect 217794 651454 218414 686898
rect 217794 650898 217826 651454
rect 218382 650898 218414 651454
rect 217794 615454 218414 650898
rect 217794 614898 217826 615454
rect 218382 614898 218414 615454
rect 217794 579454 218414 614898
rect 217794 578898 217826 579454
rect 218382 578898 218414 579454
rect 217794 543454 218414 578898
rect 217794 542898 217826 543454
rect 218382 542898 218414 543454
rect 217794 507454 218414 542898
rect 217794 506898 217826 507454
rect 218382 506898 218414 507454
rect 217794 471454 218414 506898
rect 217794 470898 217826 471454
rect 218382 470898 218414 471454
rect 217794 435454 218414 470898
rect 217794 434898 217826 435454
rect 218382 434898 218414 435454
rect 217794 399454 218414 434898
rect 217794 398898 217826 399454
rect 218382 398898 218414 399454
rect 217794 363454 218414 398898
rect 217794 362898 217826 363454
rect 218382 362898 218414 363454
rect 215888 331174 216208 331206
rect 215888 330938 215930 331174
rect 216166 330938 216208 331174
rect 215888 330854 216208 330938
rect 215888 330618 215930 330854
rect 216166 330618 216208 330854
rect 215888 330586 216208 330618
rect 207834 316938 207866 317494
rect 208422 316938 208454 317494
rect 207834 281494 208454 316938
rect 217794 327454 218414 362898
rect 217794 326898 217826 327454
rect 218382 326898 218414 327454
rect 215888 295174 216208 295206
rect 215888 294938 215930 295174
rect 216166 294938 216208 295174
rect 215888 294854 216208 294938
rect 215888 294618 215930 294854
rect 216166 294618 216208 294854
rect 215888 294586 216208 294618
rect 207834 280938 207866 281494
rect 208422 280938 208454 281494
rect 207834 245494 208454 280938
rect 217794 291454 218414 326898
rect 217794 290898 217826 291454
rect 218382 290898 218414 291454
rect 215888 259174 216208 259206
rect 215888 258938 215930 259174
rect 216166 258938 216208 259174
rect 215888 258854 216208 258938
rect 215888 258618 215930 258854
rect 216166 258618 216208 258854
rect 215888 258586 216208 258618
rect 207834 244938 207866 245494
rect 208422 244938 208454 245494
rect 207834 209494 208454 244938
rect 217794 255454 218414 290898
rect 217794 254898 217826 255454
rect 218382 254898 218414 255454
rect 215888 223174 216208 223206
rect 215888 222938 215930 223174
rect 216166 222938 216208 223174
rect 215888 222854 216208 222938
rect 215888 222618 215930 222854
rect 216166 222618 216208 222854
rect 215888 222586 216208 222618
rect 207834 208938 207866 209494
rect 208422 208938 208454 209494
rect 207834 173494 208454 208938
rect 217794 219454 218414 254898
rect 217794 218898 217826 219454
rect 218382 218898 218414 219454
rect 215888 187174 216208 187206
rect 215888 186938 215930 187174
rect 216166 186938 216208 187174
rect 215888 186854 216208 186938
rect 215888 186618 215930 186854
rect 216166 186618 216208 186854
rect 215888 186586 216208 186618
rect 207834 172938 207866 173494
rect 208422 172938 208454 173494
rect 207834 137494 208454 172938
rect 217794 183454 218414 218898
rect 217794 182898 217826 183454
rect 218382 182898 218414 183454
rect 215888 151174 216208 151206
rect 215888 150938 215930 151174
rect 216166 150938 216208 151174
rect 215888 150854 216208 150938
rect 215888 150618 215930 150854
rect 216166 150618 216208 150854
rect 215888 150586 216208 150618
rect 207834 136938 207866 137494
rect 208422 136938 208454 137494
rect 207834 101494 208454 136938
rect 217794 147454 218414 182898
rect 217794 146898 217826 147454
rect 218382 146898 218414 147454
rect 215888 115174 216208 115206
rect 215888 114938 215930 115174
rect 216166 114938 216208 115174
rect 215888 114854 216208 114938
rect 215888 114618 215930 114854
rect 216166 114618 216208 114854
rect 215888 114586 216208 114618
rect 207834 100938 207866 101494
rect 208422 100938 208454 101494
rect 207834 65494 208454 100938
rect 217794 111454 218414 146898
rect 217794 110898 217826 111454
rect 218382 110898 218414 111454
rect 215888 79174 216208 79206
rect 215888 78938 215930 79174
rect 216166 78938 216208 79174
rect 215888 78854 216208 78938
rect 215888 78618 215930 78854
rect 216166 78618 216208 78854
rect 215888 78586 216208 78618
rect 207834 64938 207866 65494
rect 208422 64938 208454 65494
rect 207834 29494 208454 64938
rect 217794 75454 218414 110898
rect 217794 74898 217826 75454
rect 218382 74898 218414 75454
rect 215888 43174 216208 43206
rect 215888 42938 215930 43174
rect 216166 42938 216208 43174
rect 215888 42854 216208 42938
rect 215888 42618 215930 42854
rect 216166 42618 216208 42854
rect 215888 42586 216208 42618
rect 207834 28938 207866 29494
rect 208422 28938 208454 29494
rect 207834 -7066 208454 28938
rect 217794 39454 218414 74898
rect 217794 38898 217826 39454
rect 218382 38898 218414 39454
rect 215888 7174 216208 7206
rect 215888 6938 215930 7174
rect 216166 6938 216208 7174
rect 215888 6854 216208 6938
rect 215888 6618 215930 6854
rect 216166 6618 216208 6854
rect 215888 6586 216208 6618
rect 207834 -7622 207866 -7066
rect 208422 -7622 208454 -7066
rect 207834 -7654 208454 -7622
rect 217794 3454 218414 38898
rect 217794 2898 217826 3454
rect 218382 2898 218414 3454
rect 217794 -346 218414 2898
rect 217794 -902 217826 -346
rect 218382 -902 218414 -346
rect 217794 -7654 218414 -902
rect 221514 705798 222134 711590
rect 221514 705242 221546 705798
rect 222102 705242 222134 705798
rect 221514 691174 222134 705242
rect 221514 690618 221546 691174
rect 222102 690618 222134 691174
rect 221514 655174 222134 690618
rect 221514 654618 221546 655174
rect 222102 654618 222134 655174
rect 221514 619174 222134 654618
rect 221514 618618 221546 619174
rect 222102 618618 222134 619174
rect 221514 583174 222134 618618
rect 221514 582618 221546 583174
rect 222102 582618 222134 583174
rect 221514 547174 222134 582618
rect 221514 546618 221546 547174
rect 222102 546618 222134 547174
rect 221514 511174 222134 546618
rect 221514 510618 221546 511174
rect 222102 510618 222134 511174
rect 221514 475174 222134 510618
rect 221514 474618 221546 475174
rect 222102 474618 222134 475174
rect 221514 439174 222134 474618
rect 221514 438618 221546 439174
rect 222102 438618 222134 439174
rect 221514 403174 222134 438618
rect 221514 402618 221546 403174
rect 222102 402618 222134 403174
rect 221514 367174 222134 402618
rect 221514 366618 221546 367174
rect 222102 366618 222134 367174
rect 221514 331174 222134 366618
rect 221514 330618 221546 331174
rect 222102 330618 222134 331174
rect 221514 295174 222134 330618
rect 221514 294618 221546 295174
rect 222102 294618 222134 295174
rect 221514 259174 222134 294618
rect 221514 258618 221546 259174
rect 222102 258618 222134 259174
rect 221514 223174 222134 258618
rect 221514 222618 221546 223174
rect 222102 222618 222134 223174
rect 221514 187174 222134 222618
rect 221514 186618 221546 187174
rect 222102 186618 222134 187174
rect 221514 151174 222134 186618
rect 221514 150618 221546 151174
rect 222102 150618 222134 151174
rect 221514 115174 222134 150618
rect 221514 114618 221546 115174
rect 222102 114618 222134 115174
rect 221514 79174 222134 114618
rect 221514 78618 221546 79174
rect 222102 78618 222134 79174
rect 221514 43174 222134 78618
rect 221514 42618 221546 43174
rect 222102 42618 222134 43174
rect 221514 7174 222134 42618
rect 221514 6618 221546 7174
rect 222102 6618 222134 7174
rect 221514 -1306 222134 6618
rect 221514 -1862 221546 -1306
rect 222102 -1862 222134 -1306
rect 221514 -7654 222134 -1862
rect 225234 706758 225854 711590
rect 225234 706202 225266 706758
rect 225822 706202 225854 706758
rect 225234 694894 225854 706202
rect 225234 694338 225266 694894
rect 225822 694338 225854 694894
rect 225234 658894 225854 694338
rect 225234 658338 225266 658894
rect 225822 658338 225854 658894
rect 225234 622894 225854 658338
rect 225234 622338 225266 622894
rect 225822 622338 225854 622894
rect 225234 586894 225854 622338
rect 225234 586338 225266 586894
rect 225822 586338 225854 586894
rect 225234 550894 225854 586338
rect 225234 550338 225266 550894
rect 225822 550338 225854 550894
rect 225234 514894 225854 550338
rect 225234 514338 225266 514894
rect 225822 514338 225854 514894
rect 225234 478894 225854 514338
rect 225234 478338 225266 478894
rect 225822 478338 225854 478894
rect 225234 442894 225854 478338
rect 225234 442338 225266 442894
rect 225822 442338 225854 442894
rect 225234 406894 225854 442338
rect 225234 406338 225266 406894
rect 225822 406338 225854 406894
rect 225234 370894 225854 406338
rect 225234 370338 225266 370894
rect 225822 370338 225854 370894
rect 225234 334894 225854 370338
rect 225234 334338 225266 334894
rect 225822 334338 225854 334894
rect 225234 298894 225854 334338
rect 225234 298338 225266 298894
rect 225822 298338 225854 298894
rect 225234 262894 225854 298338
rect 225234 262338 225266 262894
rect 225822 262338 225854 262894
rect 225234 226894 225854 262338
rect 225234 226338 225266 226894
rect 225822 226338 225854 226894
rect 225234 190894 225854 226338
rect 225234 190338 225266 190894
rect 225822 190338 225854 190894
rect 225234 154894 225854 190338
rect 225234 154338 225266 154894
rect 225822 154338 225854 154894
rect 225234 118894 225854 154338
rect 225234 118338 225266 118894
rect 225822 118338 225854 118894
rect 225234 82894 225854 118338
rect 225234 82338 225266 82894
rect 225822 82338 225854 82894
rect 225234 46894 225854 82338
rect 225234 46338 225266 46894
rect 225822 46338 225854 46894
rect 225234 10894 225854 46338
rect 225234 10338 225266 10894
rect 225822 10338 225854 10894
rect 225234 -2266 225854 10338
rect 225234 -2822 225266 -2266
rect 225822 -2822 225854 -2266
rect 225234 -7654 225854 -2822
rect 228954 707718 229574 711590
rect 228954 707162 228986 707718
rect 229542 707162 229574 707718
rect 228954 698614 229574 707162
rect 228954 698058 228986 698614
rect 229542 698058 229574 698614
rect 228954 662614 229574 698058
rect 228954 662058 228986 662614
rect 229542 662058 229574 662614
rect 228954 626614 229574 662058
rect 228954 626058 228986 626614
rect 229542 626058 229574 626614
rect 228954 590614 229574 626058
rect 228954 590058 228986 590614
rect 229542 590058 229574 590614
rect 228954 554614 229574 590058
rect 228954 554058 228986 554614
rect 229542 554058 229574 554614
rect 228954 518614 229574 554058
rect 228954 518058 228986 518614
rect 229542 518058 229574 518614
rect 228954 482614 229574 518058
rect 228954 482058 228986 482614
rect 229542 482058 229574 482614
rect 228954 446614 229574 482058
rect 228954 446058 228986 446614
rect 229542 446058 229574 446614
rect 228954 410614 229574 446058
rect 228954 410058 228986 410614
rect 229542 410058 229574 410614
rect 228954 374614 229574 410058
rect 228954 374058 228986 374614
rect 229542 374058 229574 374614
rect 228954 338614 229574 374058
rect 228954 338058 228986 338614
rect 229542 338058 229574 338614
rect 228954 302614 229574 338058
rect 232674 708678 233294 711590
rect 232674 708122 232706 708678
rect 233262 708122 233294 708678
rect 232674 666334 233294 708122
rect 232674 665778 232706 666334
rect 233262 665778 233294 666334
rect 232674 630334 233294 665778
rect 232674 629778 232706 630334
rect 233262 629778 233294 630334
rect 232674 594334 233294 629778
rect 232674 593778 232706 594334
rect 233262 593778 233294 594334
rect 232674 558334 233294 593778
rect 232674 557778 232706 558334
rect 233262 557778 233294 558334
rect 232674 522334 233294 557778
rect 232674 521778 232706 522334
rect 233262 521778 233294 522334
rect 232674 486334 233294 521778
rect 232674 485778 232706 486334
rect 233262 485778 233294 486334
rect 232674 450334 233294 485778
rect 232674 449778 232706 450334
rect 233262 449778 233294 450334
rect 232674 414334 233294 449778
rect 232674 413778 232706 414334
rect 233262 413778 233294 414334
rect 232674 378334 233294 413778
rect 232674 377778 232706 378334
rect 233262 377778 233294 378334
rect 232674 342334 233294 377778
rect 232674 341778 232706 342334
rect 233262 341778 233294 342334
rect 231248 327454 231568 327486
rect 231248 327218 231290 327454
rect 231526 327218 231568 327454
rect 231248 327134 231568 327218
rect 231248 326898 231290 327134
rect 231526 326898 231568 327134
rect 231248 326866 231568 326898
rect 228954 302058 228986 302614
rect 229542 302058 229574 302614
rect 228954 266614 229574 302058
rect 232674 306334 233294 341778
rect 232674 305778 232706 306334
rect 233262 305778 233294 306334
rect 231248 291454 231568 291486
rect 231248 291218 231290 291454
rect 231526 291218 231568 291454
rect 231248 291134 231568 291218
rect 231248 290898 231290 291134
rect 231526 290898 231568 291134
rect 231248 290866 231568 290898
rect 228954 266058 228986 266614
rect 229542 266058 229574 266614
rect 228954 230614 229574 266058
rect 232674 270334 233294 305778
rect 232674 269778 232706 270334
rect 233262 269778 233294 270334
rect 231248 255454 231568 255486
rect 231248 255218 231290 255454
rect 231526 255218 231568 255454
rect 231248 255134 231568 255218
rect 231248 254898 231290 255134
rect 231526 254898 231568 255134
rect 231248 254866 231568 254898
rect 228954 230058 228986 230614
rect 229542 230058 229574 230614
rect 228954 194614 229574 230058
rect 232674 234334 233294 269778
rect 232674 233778 232706 234334
rect 233262 233778 233294 234334
rect 231248 219454 231568 219486
rect 231248 219218 231290 219454
rect 231526 219218 231568 219454
rect 231248 219134 231568 219218
rect 231248 218898 231290 219134
rect 231526 218898 231568 219134
rect 231248 218866 231568 218898
rect 228954 194058 228986 194614
rect 229542 194058 229574 194614
rect 228954 158614 229574 194058
rect 232674 198334 233294 233778
rect 232674 197778 232706 198334
rect 233262 197778 233294 198334
rect 231248 183454 231568 183486
rect 231248 183218 231290 183454
rect 231526 183218 231568 183454
rect 231248 183134 231568 183218
rect 231248 182898 231290 183134
rect 231526 182898 231568 183134
rect 231248 182866 231568 182898
rect 228954 158058 228986 158614
rect 229542 158058 229574 158614
rect 228954 122614 229574 158058
rect 232674 162334 233294 197778
rect 232674 161778 232706 162334
rect 233262 161778 233294 162334
rect 231248 147454 231568 147486
rect 231248 147218 231290 147454
rect 231526 147218 231568 147454
rect 231248 147134 231568 147218
rect 231248 146898 231290 147134
rect 231526 146898 231568 147134
rect 231248 146866 231568 146898
rect 228954 122058 228986 122614
rect 229542 122058 229574 122614
rect 228954 86614 229574 122058
rect 232674 126334 233294 161778
rect 232674 125778 232706 126334
rect 233262 125778 233294 126334
rect 231248 111454 231568 111486
rect 231248 111218 231290 111454
rect 231526 111218 231568 111454
rect 231248 111134 231568 111218
rect 231248 110898 231290 111134
rect 231526 110898 231568 111134
rect 231248 110866 231568 110898
rect 228954 86058 228986 86614
rect 229542 86058 229574 86614
rect 228954 50614 229574 86058
rect 232674 90334 233294 125778
rect 232674 89778 232706 90334
rect 233262 89778 233294 90334
rect 231248 75454 231568 75486
rect 231248 75218 231290 75454
rect 231526 75218 231568 75454
rect 231248 75134 231568 75218
rect 231248 74898 231290 75134
rect 231526 74898 231568 75134
rect 231248 74866 231568 74898
rect 228954 50058 228986 50614
rect 229542 50058 229574 50614
rect 228954 14614 229574 50058
rect 232674 54334 233294 89778
rect 232674 53778 232706 54334
rect 233262 53778 233294 54334
rect 231248 39454 231568 39486
rect 231248 39218 231290 39454
rect 231526 39218 231568 39454
rect 231248 39134 231568 39218
rect 231248 38898 231290 39134
rect 231526 38898 231568 39134
rect 231248 38866 231568 38898
rect 228954 14058 228986 14614
rect 229542 14058 229574 14614
rect 228954 -3226 229574 14058
rect 228954 -3782 228986 -3226
rect 229542 -3782 229574 -3226
rect 228954 -7654 229574 -3782
rect 232674 18334 233294 53778
rect 232674 17778 232706 18334
rect 233262 17778 233294 18334
rect 232674 -4186 233294 17778
rect 232674 -4742 232706 -4186
rect 233262 -4742 233294 -4186
rect 232674 -7654 233294 -4742
rect 236394 709638 237014 711590
rect 236394 709082 236426 709638
rect 236982 709082 237014 709638
rect 236394 670054 237014 709082
rect 236394 669498 236426 670054
rect 236982 669498 237014 670054
rect 236394 634054 237014 669498
rect 236394 633498 236426 634054
rect 236982 633498 237014 634054
rect 236394 598054 237014 633498
rect 236394 597498 236426 598054
rect 236982 597498 237014 598054
rect 236394 562054 237014 597498
rect 236394 561498 236426 562054
rect 236982 561498 237014 562054
rect 236394 526054 237014 561498
rect 236394 525498 236426 526054
rect 236982 525498 237014 526054
rect 236394 490054 237014 525498
rect 236394 489498 236426 490054
rect 236982 489498 237014 490054
rect 236394 454054 237014 489498
rect 236394 453498 236426 454054
rect 236982 453498 237014 454054
rect 236394 418054 237014 453498
rect 236394 417498 236426 418054
rect 236982 417498 237014 418054
rect 236394 382054 237014 417498
rect 236394 381498 236426 382054
rect 236982 381498 237014 382054
rect 236394 346054 237014 381498
rect 236394 345498 236426 346054
rect 236982 345498 237014 346054
rect 236394 310054 237014 345498
rect 236394 309498 236426 310054
rect 236982 309498 237014 310054
rect 236394 274054 237014 309498
rect 236394 273498 236426 274054
rect 236982 273498 237014 274054
rect 236394 238054 237014 273498
rect 236394 237498 236426 238054
rect 236982 237498 237014 238054
rect 236394 202054 237014 237498
rect 236394 201498 236426 202054
rect 236982 201498 237014 202054
rect 236394 166054 237014 201498
rect 236394 165498 236426 166054
rect 236982 165498 237014 166054
rect 236394 130054 237014 165498
rect 236394 129498 236426 130054
rect 236982 129498 237014 130054
rect 236394 94054 237014 129498
rect 236394 93498 236426 94054
rect 236982 93498 237014 94054
rect 236394 58054 237014 93498
rect 236394 57498 236426 58054
rect 236982 57498 237014 58054
rect 236394 22054 237014 57498
rect 236394 21498 236426 22054
rect 236982 21498 237014 22054
rect 236394 -5146 237014 21498
rect 236394 -5702 236426 -5146
rect 236982 -5702 237014 -5146
rect 236394 -7654 237014 -5702
rect 240114 710598 240734 711590
rect 240114 710042 240146 710598
rect 240702 710042 240734 710598
rect 240114 673774 240734 710042
rect 240114 673218 240146 673774
rect 240702 673218 240734 673774
rect 240114 637774 240734 673218
rect 240114 637218 240146 637774
rect 240702 637218 240734 637774
rect 240114 601774 240734 637218
rect 240114 601218 240146 601774
rect 240702 601218 240734 601774
rect 240114 565774 240734 601218
rect 240114 565218 240146 565774
rect 240702 565218 240734 565774
rect 240114 529774 240734 565218
rect 240114 529218 240146 529774
rect 240702 529218 240734 529774
rect 240114 493774 240734 529218
rect 240114 493218 240146 493774
rect 240702 493218 240734 493774
rect 240114 457774 240734 493218
rect 240114 457218 240146 457774
rect 240702 457218 240734 457774
rect 240114 421774 240734 457218
rect 240114 421218 240146 421774
rect 240702 421218 240734 421774
rect 240114 385774 240734 421218
rect 240114 385218 240146 385774
rect 240702 385218 240734 385774
rect 240114 349774 240734 385218
rect 240114 349218 240146 349774
rect 240702 349218 240734 349774
rect 240114 313774 240734 349218
rect 240114 313218 240146 313774
rect 240702 313218 240734 313774
rect 240114 277774 240734 313218
rect 240114 277218 240146 277774
rect 240702 277218 240734 277774
rect 240114 241774 240734 277218
rect 240114 241218 240146 241774
rect 240702 241218 240734 241774
rect 240114 205774 240734 241218
rect 240114 205218 240146 205774
rect 240702 205218 240734 205774
rect 240114 169774 240734 205218
rect 240114 169218 240146 169774
rect 240702 169218 240734 169774
rect 240114 133774 240734 169218
rect 240114 133218 240146 133774
rect 240702 133218 240734 133774
rect 240114 97774 240734 133218
rect 240114 97218 240146 97774
rect 240702 97218 240734 97774
rect 240114 61774 240734 97218
rect 240114 61218 240146 61774
rect 240702 61218 240734 61774
rect 240114 25774 240734 61218
rect 240114 25218 240146 25774
rect 240702 25218 240734 25774
rect 240114 -6106 240734 25218
rect 240114 -6662 240146 -6106
rect 240702 -6662 240734 -6106
rect 240114 -7654 240734 -6662
rect 243834 711558 244454 711590
rect 243834 711002 243866 711558
rect 244422 711002 244454 711558
rect 243834 677494 244454 711002
rect 243834 676938 243866 677494
rect 244422 676938 244454 677494
rect 243834 641494 244454 676938
rect 243834 640938 243866 641494
rect 244422 640938 244454 641494
rect 243834 605494 244454 640938
rect 243834 604938 243866 605494
rect 244422 604938 244454 605494
rect 243834 569494 244454 604938
rect 243834 568938 243866 569494
rect 244422 568938 244454 569494
rect 243834 533494 244454 568938
rect 243834 532938 243866 533494
rect 244422 532938 244454 533494
rect 243834 497494 244454 532938
rect 243834 496938 243866 497494
rect 244422 496938 244454 497494
rect 243834 461494 244454 496938
rect 243834 460938 243866 461494
rect 244422 460938 244454 461494
rect 243834 425494 244454 460938
rect 243834 424938 243866 425494
rect 244422 424938 244454 425494
rect 243834 389494 244454 424938
rect 243834 388938 243866 389494
rect 244422 388938 244454 389494
rect 243834 353494 244454 388938
rect 243834 352938 243866 353494
rect 244422 352938 244454 353494
rect 243834 317494 244454 352938
rect 253794 704838 254414 711590
rect 253794 704282 253826 704838
rect 254382 704282 254414 704838
rect 253794 687454 254414 704282
rect 253794 686898 253826 687454
rect 254382 686898 254414 687454
rect 253794 651454 254414 686898
rect 253794 650898 253826 651454
rect 254382 650898 254414 651454
rect 253794 615454 254414 650898
rect 253794 614898 253826 615454
rect 254382 614898 254414 615454
rect 253794 579454 254414 614898
rect 253794 578898 253826 579454
rect 254382 578898 254414 579454
rect 253794 543454 254414 578898
rect 253794 542898 253826 543454
rect 254382 542898 254414 543454
rect 253794 507454 254414 542898
rect 253794 506898 253826 507454
rect 254382 506898 254414 507454
rect 253794 471454 254414 506898
rect 253794 470898 253826 471454
rect 254382 470898 254414 471454
rect 253794 435454 254414 470898
rect 253794 434898 253826 435454
rect 254382 434898 254414 435454
rect 253794 399454 254414 434898
rect 253794 398898 253826 399454
rect 254382 398898 254414 399454
rect 253794 363454 254414 398898
rect 253794 362898 253826 363454
rect 254382 362898 254414 363454
rect 246608 331174 246928 331206
rect 246608 330938 246650 331174
rect 246886 330938 246928 331174
rect 246608 330854 246928 330938
rect 246608 330618 246650 330854
rect 246886 330618 246928 330854
rect 246608 330586 246928 330618
rect 243834 316938 243866 317494
rect 244422 316938 244454 317494
rect 243834 281494 244454 316938
rect 253794 327454 254414 362898
rect 253794 326898 253826 327454
rect 254382 326898 254414 327454
rect 246608 295174 246928 295206
rect 246608 294938 246650 295174
rect 246886 294938 246928 295174
rect 246608 294854 246928 294938
rect 246608 294618 246650 294854
rect 246886 294618 246928 294854
rect 246608 294586 246928 294618
rect 243834 280938 243866 281494
rect 244422 280938 244454 281494
rect 243834 245494 244454 280938
rect 253794 291454 254414 326898
rect 253794 290898 253826 291454
rect 254382 290898 254414 291454
rect 246608 259174 246928 259206
rect 246608 258938 246650 259174
rect 246886 258938 246928 259174
rect 246608 258854 246928 258938
rect 246608 258618 246650 258854
rect 246886 258618 246928 258854
rect 246608 258586 246928 258618
rect 243834 244938 243866 245494
rect 244422 244938 244454 245494
rect 243834 209494 244454 244938
rect 253794 255454 254414 290898
rect 253794 254898 253826 255454
rect 254382 254898 254414 255454
rect 246608 223174 246928 223206
rect 246608 222938 246650 223174
rect 246886 222938 246928 223174
rect 246608 222854 246928 222938
rect 246608 222618 246650 222854
rect 246886 222618 246928 222854
rect 246608 222586 246928 222618
rect 243834 208938 243866 209494
rect 244422 208938 244454 209494
rect 243834 173494 244454 208938
rect 253794 219454 254414 254898
rect 253794 218898 253826 219454
rect 254382 218898 254414 219454
rect 246608 187174 246928 187206
rect 246608 186938 246650 187174
rect 246886 186938 246928 187174
rect 246608 186854 246928 186938
rect 246608 186618 246650 186854
rect 246886 186618 246928 186854
rect 246608 186586 246928 186618
rect 243834 172938 243866 173494
rect 244422 172938 244454 173494
rect 243834 137494 244454 172938
rect 253794 183454 254414 218898
rect 253794 182898 253826 183454
rect 254382 182898 254414 183454
rect 246608 151174 246928 151206
rect 246608 150938 246650 151174
rect 246886 150938 246928 151174
rect 246608 150854 246928 150938
rect 246608 150618 246650 150854
rect 246886 150618 246928 150854
rect 246608 150586 246928 150618
rect 243834 136938 243866 137494
rect 244422 136938 244454 137494
rect 243834 101494 244454 136938
rect 253794 147454 254414 182898
rect 253794 146898 253826 147454
rect 254382 146898 254414 147454
rect 246608 115174 246928 115206
rect 246608 114938 246650 115174
rect 246886 114938 246928 115174
rect 246608 114854 246928 114938
rect 246608 114618 246650 114854
rect 246886 114618 246928 114854
rect 246608 114586 246928 114618
rect 243834 100938 243866 101494
rect 244422 100938 244454 101494
rect 243834 65494 244454 100938
rect 253794 111454 254414 146898
rect 253794 110898 253826 111454
rect 254382 110898 254414 111454
rect 246608 79174 246928 79206
rect 246608 78938 246650 79174
rect 246886 78938 246928 79174
rect 246608 78854 246928 78938
rect 246608 78618 246650 78854
rect 246886 78618 246928 78854
rect 246608 78586 246928 78618
rect 243834 64938 243866 65494
rect 244422 64938 244454 65494
rect 243834 29494 244454 64938
rect 253794 75454 254414 110898
rect 253794 74898 253826 75454
rect 254382 74898 254414 75454
rect 246608 43174 246928 43206
rect 246608 42938 246650 43174
rect 246886 42938 246928 43174
rect 246608 42854 246928 42938
rect 246608 42618 246650 42854
rect 246886 42618 246928 42854
rect 246608 42586 246928 42618
rect 243834 28938 243866 29494
rect 244422 28938 244454 29494
rect 243834 -7066 244454 28938
rect 253794 39454 254414 74898
rect 253794 38898 253826 39454
rect 254382 38898 254414 39454
rect 246608 7174 246928 7206
rect 246608 6938 246650 7174
rect 246886 6938 246928 7174
rect 246608 6854 246928 6938
rect 246608 6618 246650 6854
rect 246886 6618 246928 6854
rect 246608 6586 246928 6618
rect 243834 -7622 243866 -7066
rect 244422 -7622 244454 -7066
rect 243834 -7654 244454 -7622
rect 253794 3454 254414 38898
rect 253794 2898 253826 3454
rect 254382 2898 254414 3454
rect 253794 -346 254414 2898
rect 253794 -902 253826 -346
rect 254382 -902 254414 -346
rect 253794 -7654 254414 -902
rect 257514 705798 258134 711590
rect 257514 705242 257546 705798
rect 258102 705242 258134 705798
rect 257514 691174 258134 705242
rect 257514 690618 257546 691174
rect 258102 690618 258134 691174
rect 257514 655174 258134 690618
rect 257514 654618 257546 655174
rect 258102 654618 258134 655174
rect 257514 619174 258134 654618
rect 257514 618618 257546 619174
rect 258102 618618 258134 619174
rect 257514 583174 258134 618618
rect 257514 582618 257546 583174
rect 258102 582618 258134 583174
rect 257514 547174 258134 582618
rect 257514 546618 257546 547174
rect 258102 546618 258134 547174
rect 257514 511174 258134 546618
rect 257514 510618 257546 511174
rect 258102 510618 258134 511174
rect 257514 475174 258134 510618
rect 257514 474618 257546 475174
rect 258102 474618 258134 475174
rect 257514 439174 258134 474618
rect 257514 438618 257546 439174
rect 258102 438618 258134 439174
rect 257514 403174 258134 438618
rect 257514 402618 257546 403174
rect 258102 402618 258134 403174
rect 257514 367174 258134 402618
rect 257514 366618 257546 367174
rect 258102 366618 258134 367174
rect 257514 331174 258134 366618
rect 261234 706758 261854 711590
rect 261234 706202 261266 706758
rect 261822 706202 261854 706758
rect 261234 694894 261854 706202
rect 261234 694338 261266 694894
rect 261822 694338 261854 694894
rect 261234 658894 261854 694338
rect 261234 658338 261266 658894
rect 261822 658338 261854 658894
rect 261234 622894 261854 658338
rect 261234 622338 261266 622894
rect 261822 622338 261854 622894
rect 261234 586894 261854 622338
rect 261234 586338 261266 586894
rect 261822 586338 261854 586894
rect 261234 550894 261854 586338
rect 261234 550338 261266 550894
rect 261822 550338 261854 550894
rect 261234 514894 261854 550338
rect 261234 514338 261266 514894
rect 261822 514338 261854 514894
rect 261234 478894 261854 514338
rect 261234 478338 261266 478894
rect 261822 478338 261854 478894
rect 261234 442894 261854 478338
rect 261234 442338 261266 442894
rect 261822 442338 261854 442894
rect 261234 406894 261854 442338
rect 261234 406338 261266 406894
rect 261822 406338 261854 406894
rect 261234 370894 261854 406338
rect 261234 370338 261266 370894
rect 261822 370338 261854 370894
rect 261234 354980 261854 370338
rect 264954 707718 265574 711590
rect 264954 707162 264986 707718
rect 265542 707162 265574 707718
rect 264954 698614 265574 707162
rect 264954 698058 264986 698614
rect 265542 698058 265574 698614
rect 264954 662614 265574 698058
rect 264954 662058 264986 662614
rect 265542 662058 265574 662614
rect 264954 626614 265574 662058
rect 264954 626058 264986 626614
rect 265542 626058 265574 626614
rect 264954 590614 265574 626058
rect 264954 590058 264986 590614
rect 265542 590058 265574 590614
rect 264954 554614 265574 590058
rect 264954 554058 264986 554614
rect 265542 554058 265574 554614
rect 264954 518614 265574 554058
rect 264954 518058 264986 518614
rect 265542 518058 265574 518614
rect 264954 482614 265574 518058
rect 264954 482058 264986 482614
rect 265542 482058 265574 482614
rect 264954 446614 265574 482058
rect 264954 446058 264986 446614
rect 265542 446058 265574 446614
rect 264954 410614 265574 446058
rect 264954 410058 264986 410614
rect 265542 410058 265574 410614
rect 264954 374614 265574 410058
rect 264954 374058 264986 374614
rect 265542 374058 265574 374614
rect 257514 330618 257546 331174
rect 258102 330618 258134 331174
rect 257514 295174 258134 330618
rect 264954 338614 265574 374058
rect 264954 338058 264986 338614
rect 265542 338058 265574 338614
rect 261968 327454 262288 327486
rect 261968 327218 262010 327454
rect 262246 327218 262288 327454
rect 261968 327134 262288 327218
rect 261968 326898 262010 327134
rect 262246 326898 262288 327134
rect 261968 326866 262288 326898
rect 257514 294618 257546 295174
rect 258102 294618 258134 295174
rect 257514 259174 258134 294618
rect 264954 302614 265574 338058
rect 264954 302058 264986 302614
rect 265542 302058 265574 302614
rect 261968 291454 262288 291486
rect 261968 291218 262010 291454
rect 262246 291218 262288 291454
rect 261968 291134 262288 291218
rect 261968 290898 262010 291134
rect 262246 290898 262288 291134
rect 261968 290866 262288 290898
rect 257514 258618 257546 259174
rect 258102 258618 258134 259174
rect 257514 223174 258134 258618
rect 264954 266614 265574 302058
rect 264954 266058 264986 266614
rect 265542 266058 265574 266614
rect 261968 255454 262288 255486
rect 261968 255218 262010 255454
rect 262246 255218 262288 255454
rect 261968 255134 262288 255218
rect 261968 254898 262010 255134
rect 262246 254898 262288 255134
rect 261968 254866 262288 254898
rect 257514 222618 257546 223174
rect 258102 222618 258134 223174
rect 257514 187174 258134 222618
rect 264954 230614 265574 266058
rect 264954 230058 264986 230614
rect 265542 230058 265574 230614
rect 261968 219454 262288 219486
rect 261968 219218 262010 219454
rect 262246 219218 262288 219454
rect 261968 219134 262288 219218
rect 261968 218898 262010 219134
rect 262246 218898 262288 219134
rect 261968 218866 262288 218898
rect 257514 186618 257546 187174
rect 258102 186618 258134 187174
rect 257514 151174 258134 186618
rect 264954 194614 265574 230058
rect 264954 194058 264986 194614
rect 265542 194058 265574 194614
rect 261968 183454 262288 183486
rect 261968 183218 262010 183454
rect 262246 183218 262288 183454
rect 261968 183134 262288 183218
rect 261968 182898 262010 183134
rect 262246 182898 262288 183134
rect 261968 182866 262288 182898
rect 257514 150618 257546 151174
rect 258102 150618 258134 151174
rect 257514 115174 258134 150618
rect 264954 158614 265574 194058
rect 264954 158058 264986 158614
rect 265542 158058 265574 158614
rect 261968 147454 262288 147486
rect 261968 147218 262010 147454
rect 262246 147218 262288 147454
rect 261968 147134 262288 147218
rect 261968 146898 262010 147134
rect 262246 146898 262288 147134
rect 261968 146866 262288 146898
rect 257514 114618 257546 115174
rect 258102 114618 258134 115174
rect 257514 79174 258134 114618
rect 264954 122614 265574 158058
rect 264954 122058 264986 122614
rect 265542 122058 265574 122614
rect 261968 111454 262288 111486
rect 261968 111218 262010 111454
rect 262246 111218 262288 111454
rect 261968 111134 262288 111218
rect 261968 110898 262010 111134
rect 262246 110898 262288 111134
rect 261968 110866 262288 110898
rect 257514 78618 257546 79174
rect 258102 78618 258134 79174
rect 257514 43174 258134 78618
rect 264954 86614 265574 122058
rect 264954 86058 264986 86614
rect 265542 86058 265574 86614
rect 261968 75454 262288 75486
rect 261968 75218 262010 75454
rect 262246 75218 262288 75454
rect 261968 75134 262288 75218
rect 261968 74898 262010 75134
rect 262246 74898 262288 75134
rect 261968 74866 262288 74898
rect 257514 42618 257546 43174
rect 258102 42618 258134 43174
rect 257514 7174 258134 42618
rect 264954 50614 265574 86058
rect 264954 50058 264986 50614
rect 265542 50058 265574 50614
rect 261968 39454 262288 39486
rect 261968 39218 262010 39454
rect 262246 39218 262288 39454
rect 261968 39134 262288 39218
rect 261968 38898 262010 39134
rect 262246 38898 262288 39134
rect 261968 38866 262288 38898
rect 257514 6618 257546 7174
rect 258102 6618 258134 7174
rect 257514 -1306 258134 6618
rect 257514 -1862 257546 -1306
rect 258102 -1862 258134 -1306
rect 257514 -7654 258134 -1862
rect 264954 14614 265574 50058
rect 264954 14058 264986 14614
rect 265542 14058 265574 14614
rect 264954 -3226 265574 14058
rect 264954 -3782 264986 -3226
rect 265542 -3782 265574 -3226
rect 264954 -7654 265574 -3782
rect 268674 708678 269294 711590
rect 268674 708122 268706 708678
rect 269262 708122 269294 708678
rect 268674 666334 269294 708122
rect 268674 665778 268706 666334
rect 269262 665778 269294 666334
rect 268674 630334 269294 665778
rect 268674 629778 268706 630334
rect 269262 629778 269294 630334
rect 268674 594334 269294 629778
rect 268674 593778 268706 594334
rect 269262 593778 269294 594334
rect 268674 558334 269294 593778
rect 268674 557778 268706 558334
rect 269262 557778 269294 558334
rect 268674 522334 269294 557778
rect 268674 521778 268706 522334
rect 269262 521778 269294 522334
rect 268674 486334 269294 521778
rect 268674 485778 268706 486334
rect 269262 485778 269294 486334
rect 268674 450334 269294 485778
rect 268674 449778 268706 450334
rect 269262 449778 269294 450334
rect 268674 414334 269294 449778
rect 268674 413778 268706 414334
rect 269262 413778 269294 414334
rect 268674 378334 269294 413778
rect 268674 377778 268706 378334
rect 269262 377778 269294 378334
rect 268674 342334 269294 377778
rect 268674 341778 268706 342334
rect 269262 341778 269294 342334
rect 268674 306334 269294 341778
rect 268674 305778 268706 306334
rect 269262 305778 269294 306334
rect 268674 270334 269294 305778
rect 268674 269778 268706 270334
rect 269262 269778 269294 270334
rect 268674 234334 269294 269778
rect 268674 233778 268706 234334
rect 269262 233778 269294 234334
rect 268674 198334 269294 233778
rect 268674 197778 268706 198334
rect 269262 197778 269294 198334
rect 268674 162334 269294 197778
rect 268674 161778 268706 162334
rect 269262 161778 269294 162334
rect 268674 126334 269294 161778
rect 268674 125778 268706 126334
rect 269262 125778 269294 126334
rect 268674 90334 269294 125778
rect 268674 89778 268706 90334
rect 269262 89778 269294 90334
rect 268674 54334 269294 89778
rect 268674 53778 268706 54334
rect 269262 53778 269294 54334
rect 268674 18334 269294 53778
rect 268674 17778 268706 18334
rect 269262 17778 269294 18334
rect 268674 -4186 269294 17778
rect 268674 -4742 268706 -4186
rect 269262 -4742 269294 -4186
rect 268674 -7654 269294 -4742
rect 272394 709638 273014 711590
rect 272394 709082 272426 709638
rect 272982 709082 273014 709638
rect 272394 670054 273014 709082
rect 272394 669498 272426 670054
rect 272982 669498 273014 670054
rect 272394 634054 273014 669498
rect 272394 633498 272426 634054
rect 272982 633498 273014 634054
rect 272394 598054 273014 633498
rect 272394 597498 272426 598054
rect 272982 597498 273014 598054
rect 272394 562054 273014 597498
rect 272394 561498 272426 562054
rect 272982 561498 273014 562054
rect 272394 526054 273014 561498
rect 272394 525498 272426 526054
rect 272982 525498 273014 526054
rect 272394 490054 273014 525498
rect 272394 489498 272426 490054
rect 272982 489498 273014 490054
rect 272394 454054 273014 489498
rect 272394 453498 272426 454054
rect 272982 453498 273014 454054
rect 272394 418054 273014 453498
rect 272394 417498 272426 418054
rect 272982 417498 273014 418054
rect 272394 382054 273014 417498
rect 272394 381498 272426 382054
rect 272982 381498 273014 382054
rect 272394 346054 273014 381498
rect 272394 345498 272426 346054
rect 272982 345498 273014 346054
rect 272394 310054 273014 345498
rect 272394 309498 272426 310054
rect 272982 309498 273014 310054
rect 272394 274054 273014 309498
rect 272394 273498 272426 274054
rect 272982 273498 273014 274054
rect 272394 238054 273014 273498
rect 272394 237498 272426 238054
rect 272982 237498 273014 238054
rect 272394 202054 273014 237498
rect 272394 201498 272426 202054
rect 272982 201498 273014 202054
rect 272394 166054 273014 201498
rect 272394 165498 272426 166054
rect 272982 165498 273014 166054
rect 272394 130054 273014 165498
rect 272394 129498 272426 130054
rect 272982 129498 273014 130054
rect 272394 94054 273014 129498
rect 272394 93498 272426 94054
rect 272982 93498 273014 94054
rect 272394 58054 273014 93498
rect 272394 57498 272426 58054
rect 272982 57498 273014 58054
rect 272394 22054 273014 57498
rect 272394 21498 272426 22054
rect 272982 21498 273014 22054
rect 272394 -5146 273014 21498
rect 272394 -5702 272426 -5146
rect 272982 -5702 273014 -5146
rect 272394 -7654 273014 -5702
rect 276114 710598 276734 711590
rect 276114 710042 276146 710598
rect 276702 710042 276734 710598
rect 276114 673774 276734 710042
rect 276114 673218 276146 673774
rect 276702 673218 276734 673774
rect 276114 637774 276734 673218
rect 276114 637218 276146 637774
rect 276702 637218 276734 637774
rect 276114 601774 276734 637218
rect 276114 601218 276146 601774
rect 276702 601218 276734 601774
rect 276114 565774 276734 601218
rect 276114 565218 276146 565774
rect 276702 565218 276734 565774
rect 276114 529774 276734 565218
rect 276114 529218 276146 529774
rect 276702 529218 276734 529774
rect 276114 493774 276734 529218
rect 276114 493218 276146 493774
rect 276702 493218 276734 493774
rect 276114 457774 276734 493218
rect 276114 457218 276146 457774
rect 276702 457218 276734 457774
rect 276114 421774 276734 457218
rect 276114 421218 276146 421774
rect 276702 421218 276734 421774
rect 276114 385774 276734 421218
rect 276114 385218 276146 385774
rect 276702 385218 276734 385774
rect 276114 349774 276734 385218
rect 276114 349218 276146 349774
rect 276702 349218 276734 349774
rect 276114 313774 276734 349218
rect 279834 711558 280454 711590
rect 279834 711002 279866 711558
rect 280422 711002 280454 711558
rect 279834 677494 280454 711002
rect 279834 676938 279866 677494
rect 280422 676938 280454 677494
rect 279834 641494 280454 676938
rect 279834 640938 279866 641494
rect 280422 640938 280454 641494
rect 279834 605494 280454 640938
rect 279834 604938 279866 605494
rect 280422 604938 280454 605494
rect 279834 569494 280454 604938
rect 279834 568938 279866 569494
rect 280422 568938 280454 569494
rect 279834 533494 280454 568938
rect 279834 532938 279866 533494
rect 280422 532938 280454 533494
rect 279834 497494 280454 532938
rect 279834 496938 279866 497494
rect 280422 496938 280454 497494
rect 279834 461494 280454 496938
rect 279834 460938 279866 461494
rect 280422 460938 280454 461494
rect 279834 425494 280454 460938
rect 279834 424938 279866 425494
rect 280422 424938 280454 425494
rect 279834 389494 280454 424938
rect 279834 388938 279866 389494
rect 280422 388938 280454 389494
rect 279834 353494 280454 388938
rect 279834 352938 279866 353494
rect 280422 352938 280454 353494
rect 277328 331174 277648 331206
rect 277328 330938 277370 331174
rect 277606 330938 277648 331174
rect 277328 330854 277648 330938
rect 277328 330618 277370 330854
rect 277606 330618 277648 330854
rect 277328 330586 277648 330618
rect 276114 313218 276146 313774
rect 276702 313218 276734 313774
rect 276114 277774 276734 313218
rect 279834 317494 280454 352938
rect 279834 316938 279866 317494
rect 280422 316938 280454 317494
rect 277328 295174 277648 295206
rect 277328 294938 277370 295174
rect 277606 294938 277648 295174
rect 277328 294854 277648 294938
rect 277328 294618 277370 294854
rect 277606 294618 277648 294854
rect 277328 294586 277648 294618
rect 276114 277218 276146 277774
rect 276702 277218 276734 277774
rect 276114 241774 276734 277218
rect 279834 281494 280454 316938
rect 279834 280938 279866 281494
rect 280422 280938 280454 281494
rect 277328 259174 277648 259206
rect 277328 258938 277370 259174
rect 277606 258938 277648 259174
rect 277328 258854 277648 258938
rect 277328 258618 277370 258854
rect 277606 258618 277648 258854
rect 277328 258586 277648 258618
rect 276114 241218 276146 241774
rect 276702 241218 276734 241774
rect 276114 205774 276734 241218
rect 279834 245494 280454 280938
rect 279834 244938 279866 245494
rect 280422 244938 280454 245494
rect 277328 223174 277648 223206
rect 277328 222938 277370 223174
rect 277606 222938 277648 223174
rect 277328 222854 277648 222938
rect 277328 222618 277370 222854
rect 277606 222618 277648 222854
rect 277328 222586 277648 222618
rect 276114 205218 276146 205774
rect 276702 205218 276734 205774
rect 276114 169774 276734 205218
rect 279834 209494 280454 244938
rect 279834 208938 279866 209494
rect 280422 208938 280454 209494
rect 277328 187174 277648 187206
rect 277328 186938 277370 187174
rect 277606 186938 277648 187174
rect 277328 186854 277648 186938
rect 277328 186618 277370 186854
rect 277606 186618 277648 186854
rect 277328 186586 277648 186618
rect 276114 169218 276146 169774
rect 276702 169218 276734 169774
rect 276114 133774 276734 169218
rect 279834 173494 280454 208938
rect 279834 172938 279866 173494
rect 280422 172938 280454 173494
rect 277328 151174 277648 151206
rect 277328 150938 277370 151174
rect 277606 150938 277648 151174
rect 277328 150854 277648 150938
rect 277328 150618 277370 150854
rect 277606 150618 277648 150854
rect 277328 150586 277648 150618
rect 276114 133218 276146 133774
rect 276702 133218 276734 133774
rect 276114 97774 276734 133218
rect 279834 137494 280454 172938
rect 279834 136938 279866 137494
rect 280422 136938 280454 137494
rect 277328 115174 277648 115206
rect 277328 114938 277370 115174
rect 277606 114938 277648 115174
rect 277328 114854 277648 114938
rect 277328 114618 277370 114854
rect 277606 114618 277648 114854
rect 277328 114586 277648 114618
rect 276114 97218 276146 97774
rect 276702 97218 276734 97774
rect 276114 61774 276734 97218
rect 279834 101494 280454 136938
rect 279834 100938 279866 101494
rect 280422 100938 280454 101494
rect 277328 79174 277648 79206
rect 277328 78938 277370 79174
rect 277606 78938 277648 79174
rect 277328 78854 277648 78938
rect 277328 78618 277370 78854
rect 277606 78618 277648 78854
rect 277328 78586 277648 78618
rect 276114 61218 276146 61774
rect 276702 61218 276734 61774
rect 276114 25774 276734 61218
rect 279834 65494 280454 100938
rect 279834 64938 279866 65494
rect 280422 64938 280454 65494
rect 277328 43174 277648 43206
rect 277328 42938 277370 43174
rect 277606 42938 277648 43174
rect 277328 42854 277648 42938
rect 277328 42618 277370 42854
rect 277606 42618 277648 42854
rect 277328 42586 277648 42618
rect 276114 25218 276146 25774
rect 276702 25218 276734 25774
rect 276114 -6106 276734 25218
rect 279834 29494 280454 64938
rect 279834 28938 279866 29494
rect 280422 28938 280454 29494
rect 277328 7174 277648 7206
rect 277328 6938 277370 7174
rect 277606 6938 277648 7174
rect 277328 6854 277648 6938
rect 277328 6618 277370 6854
rect 277606 6618 277648 6854
rect 277328 6586 277648 6618
rect 276114 -6662 276146 -6106
rect 276702 -6662 276734 -6106
rect 276114 -7654 276734 -6662
rect 279834 -7066 280454 28938
rect 279834 -7622 279866 -7066
rect 280422 -7622 280454 -7066
rect 279834 -7654 280454 -7622
rect 289794 704838 290414 711590
rect 289794 704282 289826 704838
rect 290382 704282 290414 704838
rect 289794 687454 290414 704282
rect 289794 686898 289826 687454
rect 290382 686898 290414 687454
rect 289794 651454 290414 686898
rect 289794 650898 289826 651454
rect 290382 650898 290414 651454
rect 289794 615454 290414 650898
rect 289794 614898 289826 615454
rect 290382 614898 290414 615454
rect 289794 579454 290414 614898
rect 289794 578898 289826 579454
rect 290382 578898 290414 579454
rect 289794 543454 290414 578898
rect 289794 542898 289826 543454
rect 290382 542898 290414 543454
rect 289794 507454 290414 542898
rect 289794 506898 289826 507454
rect 290382 506898 290414 507454
rect 289794 471454 290414 506898
rect 289794 470898 289826 471454
rect 290382 470898 290414 471454
rect 289794 435454 290414 470898
rect 289794 434898 289826 435454
rect 290382 434898 290414 435454
rect 289794 399454 290414 434898
rect 289794 398898 289826 399454
rect 290382 398898 290414 399454
rect 289794 363454 290414 398898
rect 289794 362898 289826 363454
rect 290382 362898 290414 363454
rect 289794 327454 290414 362898
rect 293514 705798 294134 711590
rect 293514 705242 293546 705798
rect 294102 705242 294134 705798
rect 293514 691174 294134 705242
rect 293514 690618 293546 691174
rect 294102 690618 294134 691174
rect 293514 655174 294134 690618
rect 293514 654618 293546 655174
rect 294102 654618 294134 655174
rect 293514 619174 294134 654618
rect 293514 618618 293546 619174
rect 294102 618618 294134 619174
rect 293514 583174 294134 618618
rect 293514 582618 293546 583174
rect 294102 582618 294134 583174
rect 293514 547174 294134 582618
rect 293514 546618 293546 547174
rect 294102 546618 294134 547174
rect 293514 511174 294134 546618
rect 293514 510618 293546 511174
rect 294102 510618 294134 511174
rect 293514 475174 294134 510618
rect 293514 474618 293546 475174
rect 294102 474618 294134 475174
rect 293514 439174 294134 474618
rect 293514 438618 293546 439174
rect 294102 438618 294134 439174
rect 293514 403174 294134 438618
rect 293514 402618 293546 403174
rect 294102 402618 294134 403174
rect 293514 367174 294134 402618
rect 293514 366618 293546 367174
rect 294102 366618 294134 367174
rect 293514 331174 294134 366618
rect 293514 330618 293546 331174
rect 294102 330618 294134 331174
rect 289794 326898 289826 327454
rect 290382 326898 290414 327454
rect 289794 291454 290414 326898
rect 292688 327454 293008 327486
rect 292688 327218 292730 327454
rect 292966 327218 293008 327454
rect 292688 327134 293008 327218
rect 292688 326898 292730 327134
rect 292966 326898 293008 327134
rect 292688 326866 293008 326898
rect 293514 295174 294134 330618
rect 293514 294618 293546 295174
rect 294102 294618 294134 295174
rect 289794 290898 289826 291454
rect 290382 290898 290414 291454
rect 289794 255454 290414 290898
rect 292688 291454 293008 291486
rect 292688 291218 292730 291454
rect 292966 291218 293008 291454
rect 292688 291134 293008 291218
rect 292688 290898 292730 291134
rect 292966 290898 293008 291134
rect 292688 290866 293008 290898
rect 293514 259174 294134 294618
rect 293514 258618 293546 259174
rect 294102 258618 294134 259174
rect 289794 254898 289826 255454
rect 290382 254898 290414 255454
rect 289794 219454 290414 254898
rect 292688 255454 293008 255486
rect 292688 255218 292730 255454
rect 292966 255218 293008 255454
rect 292688 255134 293008 255218
rect 292688 254898 292730 255134
rect 292966 254898 293008 255134
rect 292688 254866 293008 254898
rect 293514 223174 294134 258618
rect 293514 222618 293546 223174
rect 294102 222618 294134 223174
rect 289794 218898 289826 219454
rect 290382 218898 290414 219454
rect 289794 183454 290414 218898
rect 292688 219454 293008 219486
rect 292688 219218 292730 219454
rect 292966 219218 293008 219454
rect 292688 219134 293008 219218
rect 292688 218898 292730 219134
rect 292966 218898 293008 219134
rect 292688 218866 293008 218898
rect 293514 187174 294134 222618
rect 293514 186618 293546 187174
rect 294102 186618 294134 187174
rect 289794 182898 289826 183454
rect 290382 182898 290414 183454
rect 289794 147454 290414 182898
rect 292688 183454 293008 183486
rect 292688 183218 292730 183454
rect 292966 183218 293008 183454
rect 292688 183134 293008 183218
rect 292688 182898 292730 183134
rect 292966 182898 293008 183134
rect 292688 182866 293008 182898
rect 293514 151174 294134 186618
rect 293514 150618 293546 151174
rect 294102 150618 294134 151174
rect 289794 146898 289826 147454
rect 290382 146898 290414 147454
rect 289794 111454 290414 146898
rect 292688 147454 293008 147486
rect 292688 147218 292730 147454
rect 292966 147218 293008 147454
rect 292688 147134 293008 147218
rect 292688 146898 292730 147134
rect 292966 146898 293008 147134
rect 292688 146866 293008 146898
rect 293514 115174 294134 150618
rect 293514 114618 293546 115174
rect 294102 114618 294134 115174
rect 289794 110898 289826 111454
rect 290382 110898 290414 111454
rect 289794 75454 290414 110898
rect 292688 111454 293008 111486
rect 292688 111218 292730 111454
rect 292966 111218 293008 111454
rect 292688 111134 293008 111218
rect 292688 110898 292730 111134
rect 292966 110898 293008 111134
rect 292688 110866 293008 110898
rect 293514 79174 294134 114618
rect 293514 78618 293546 79174
rect 294102 78618 294134 79174
rect 289794 74898 289826 75454
rect 290382 74898 290414 75454
rect 289794 39454 290414 74898
rect 292688 75454 293008 75486
rect 292688 75218 292730 75454
rect 292966 75218 293008 75454
rect 292688 75134 293008 75218
rect 292688 74898 292730 75134
rect 292966 74898 293008 75134
rect 292688 74866 293008 74898
rect 293514 43174 294134 78618
rect 293514 42618 293546 43174
rect 294102 42618 294134 43174
rect 289794 38898 289826 39454
rect 290382 38898 290414 39454
rect 289794 3454 290414 38898
rect 292688 39454 293008 39486
rect 292688 39218 292730 39454
rect 292966 39218 293008 39454
rect 292688 39134 293008 39218
rect 292688 38898 292730 39134
rect 292966 38898 293008 39134
rect 292688 38866 293008 38898
rect 289794 2898 289826 3454
rect 290382 2898 290414 3454
rect 289794 -346 290414 2898
rect 289794 -902 289826 -346
rect 290382 -902 290414 -346
rect 289794 -7654 290414 -902
rect 293514 7174 294134 42618
rect 293514 6618 293546 7174
rect 294102 6618 294134 7174
rect 293514 -1306 294134 6618
rect 293514 -1862 293546 -1306
rect 294102 -1862 294134 -1306
rect 293514 -7654 294134 -1862
rect 297234 706758 297854 711590
rect 297234 706202 297266 706758
rect 297822 706202 297854 706758
rect 297234 694894 297854 706202
rect 297234 694338 297266 694894
rect 297822 694338 297854 694894
rect 297234 658894 297854 694338
rect 297234 658338 297266 658894
rect 297822 658338 297854 658894
rect 297234 622894 297854 658338
rect 297234 622338 297266 622894
rect 297822 622338 297854 622894
rect 297234 586894 297854 622338
rect 297234 586338 297266 586894
rect 297822 586338 297854 586894
rect 297234 550894 297854 586338
rect 297234 550338 297266 550894
rect 297822 550338 297854 550894
rect 297234 514894 297854 550338
rect 297234 514338 297266 514894
rect 297822 514338 297854 514894
rect 297234 478894 297854 514338
rect 297234 478338 297266 478894
rect 297822 478338 297854 478894
rect 297234 442894 297854 478338
rect 297234 442338 297266 442894
rect 297822 442338 297854 442894
rect 297234 406894 297854 442338
rect 297234 406338 297266 406894
rect 297822 406338 297854 406894
rect 297234 370894 297854 406338
rect 297234 370338 297266 370894
rect 297822 370338 297854 370894
rect 297234 334894 297854 370338
rect 297234 334338 297266 334894
rect 297822 334338 297854 334894
rect 297234 298894 297854 334338
rect 297234 298338 297266 298894
rect 297822 298338 297854 298894
rect 297234 262894 297854 298338
rect 297234 262338 297266 262894
rect 297822 262338 297854 262894
rect 297234 226894 297854 262338
rect 297234 226338 297266 226894
rect 297822 226338 297854 226894
rect 297234 190894 297854 226338
rect 297234 190338 297266 190894
rect 297822 190338 297854 190894
rect 297234 154894 297854 190338
rect 297234 154338 297266 154894
rect 297822 154338 297854 154894
rect 297234 118894 297854 154338
rect 297234 118338 297266 118894
rect 297822 118338 297854 118894
rect 297234 82894 297854 118338
rect 297234 82338 297266 82894
rect 297822 82338 297854 82894
rect 297234 46894 297854 82338
rect 297234 46338 297266 46894
rect 297822 46338 297854 46894
rect 297234 10894 297854 46338
rect 297234 10338 297266 10894
rect 297822 10338 297854 10894
rect 297234 -2266 297854 10338
rect 297234 -2822 297266 -2266
rect 297822 -2822 297854 -2266
rect 297234 -7654 297854 -2822
rect 300954 707718 301574 711590
rect 300954 707162 300986 707718
rect 301542 707162 301574 707718
rect 300954 698614 301574 707162
rect 300954 698058 300986 698614
rect 301542 698058 301574 698614
rect 300954 662614 301574 698058
rect 300954 662058 300986 662614
rect 301542 662058 301574 662614
rect 300954 626614 301574 662058
rect 300954 626058 300986 626614
rect 301542 626058 301574 626614
rect 300954 590614 301574 626058
rect 300954 590058 300986 590614
rect 301542 590058 301574 590614
rect 300954 554614 301574 590058
rect 300954 554058 300986 554614
rect 301542 554058 301574 554614
rect 300954 518614 301574 554058
rect 300954 518058 300986 518614
rect 301542 518058 301574 518614
rect 300954 482614 301574 518058
rect 300954 482058 300986 482614
rect 301542 482058 301574 482614
rect 300954 446614 301574 482058
rect 300954 446058 300986 446614
rect 301542 446058 301574 446614
rect 300954 410614 301574 446058
rect 300954 410058 300986 410614
rect 301542 410058 301574 410614
rect 300954 374614 301574 410058
rect 300954 374058 300986 374614
rect 301542 374058 301574 374614
rect 300954 338614 301574 374058
rect 300954 338058 300986 338614
rect 301542 338058 301574 338614
rect 300954 302614 301574 338058
rect 300954 302058 300986 302614
rect 301542 302058 301574 302614
rect 300954 266614 301574 302058
rect 300954 266058 300986 266614
rect 301542 266058 301574 266614
rect 300954 230614 301574 266058
rect 300954 230058 300986 230614
rect 301542 230058 301574 230614
rect 300954 194614 301574 230058
rect 300954 194058 300986 194614
rect 301542 194058 301574 194614
rect 300954 158614 301574 194058
rect 300954 158058 300986 158614
rect 301542 158058 301574 158614
rect 300954 122614 301574 158058
rect 300954 122058 300986 122614
rect 301542 122058 301574 122614
rect 300954 86614 301574 122058
rect 300954 86058 300986 86614
rect 301542 86058 301574 86614
rect 300954 50614 301574 86058
rect 300954 50058 300986 50614
rect 301542 50058 301574 50614
rect 300954 14614 301574 50058
rect 300954 14058 300986 14614
rect 301542 14058 301574 14614
rect 300954 -3226 301574 14058
rect 300954 -3782 300986 -3226
rect 301542 -3782 301574 -3226
rect 300954 -7654 301574 -3782
rect 304674 708678 305294 711590
rect 304674 708122 304706 708678
rect 305262 708122 305294 708678
rect 304674 666334 305294 708122
rect 304674 665778 304706 666334
rect 305262 665778 305294 666334
rect 304674 630334 305294 665778
rect 304674 629778 304706 630334
rect 305262 629778 305294 630334
rect 304674 594334 305294 629778
rect 304674 593778 304706 594334
rect 305262 593778 305294 594334
rect 304674 558334 305294 593778
rect 304674 557778 304706 558334
rect 305262 557778 305294 558334
rect 304674 522334 305294 557778
rect 304674 521778 304706 522334
rect 305262 521778 305294 522334
rect 304674 486334 305294 521778
rect 304674 485778 304706 486334
rect 305262 485778 305294 486334
rect 304674 450334 305294 485778
rect 304674 449778 304706 450334
rect 305262 449778 305294 450334
rect 304674 414334 305294 449778
rect 304674 413778 304706 414334
rect 305262 413778 305294 414334
rect 304674 378334 305294 413778
rect 304674 377778 304706 378334
rect 305262 377778 305294 378334
rect 304674 342334 305294 377778
rect 308394 709638 309014 711590
rect 308394 709082 308426 709638
rect 308982 709082 309014 709638
rect 308394 670054 309014 709082
rect 308394 669498 308426 670054
rect 308982 669498 309014 670054
rect 308394 634054 309014 669498
rect 308394 633498 308426 634054
rect 308982 633498 309014 634054
rect 308394 598054 309014 633498
rect 308394 597498 308426 598054
rect 308982 597498 309014 598054
rect 308394 562054 309014 597498
rect 308394 561498 308426 562054
rect 308982 561498 309014 562054
rect 308394 526054 309014 561498
rect 308394 525498 308426 526054
rect 308982 525498 309014 526054
rect 308394 490054 309014 525498
rect 308394 489498 308426 490054
rect 308982 489498 309014 490054
rect 308394 454054 309014 489498
rect 308394 453498 308426 454054
rect 308982 453498 309014 454054
rect 308394 418054 309014 453498
rect 308394 417498 308426 418054
rect 308982 417498 309014 418054
rect 308394 382054 309014 417498
rect 308394 381498 308426 382054
rect 308982 381498 309014 382054
rect 308394 354980 309014 381498
rect 312114 710598 312734 711590
rect 312114 710042 312146 710598
rect 312702 710042 312734 710598
rect 312114 673774 312734 710042
rect 312114 673218 312146 673774
rect 312702 673218 312734 673774
rect 312114 637774 312734 673218
rect 312114 637218 312146 637774
rect 312702 637218 312734 637774
rect 312114 601774 312734 637218
rect 312114 601218 312146 601774
rect 312702 601218 312734 601774
rect 312114 565774 312734 601218
rect 312114 565218 312146 565774
rect 312702 565218 312734 565774
rect 312114 529774 312734 565218
rect 312114 529218 312146 529774
rect 312702 529218 312734 529774
rect 312114 493774 312734 529218
rect 312114 493218 312146 493774
rect 312702 493218 312734 493774
rect 312114 457774 312734 493218
rect 312114 457218 312146 457774
rect 312702 457218 312734 457774
rect 312114 421774 312734 457218
rect 312114 421218 312146 421774
rect 312702 421218 312734 421774
rect 312114 385774 312734 421218
rect 312114 385218 312146 385774
rect 312702 385218 312734 385774
rect 304674 341778 304706 342334
rect 305262 341778 305294 342334
rect 304674 306334 305294 341778
rect 312114 349774 312734 385218
rect 312114 349218 312146 349774
rect 312702 349218 312734 349774
rect 308048 331174 308368 331206
rect 308048 330938 308090 331174
rect 308326 330938 308368 331174
rect 308048 330854 308368 330938
rect 308048 330618 308090 330854
rect 308326 330618 308368 330854
rect 308048 330586 308368 330618
rect 304674 305778 304706 306334
rect 305262 305778 305294 306334
rect 304674 270334 305294 305778
rect 312114 313774 312734 349218
rect 312114 313218 312146 313774
rect 312702 313218 312734 313774
rect 308048 295174 308368 295206
rect 308048 294938 308090 295174
rect 308326 294938 308368 295174
rect 308048 294854 308368 294938
rect 308048 294618 308090 294854
rect 308326 294618 308368 294854
rect 308048 294586 308368 294618
rect 304674 269778 304706 270334
rect 305262 269778 305294 270334
rect 304674 234334 305294 269778
rect 312114 277774 312734 313218
rect 312114 277218 312146 277774
rect 312702 277218 312734 277774
rect 308048 259174 308368 259206
rect 308048 258938 308090 259174
rect 308326 258938 308368 259174
rect 308048 258854 308368 258938
rect 308048 258618 308090 258854
rect 308326 258618 308368 258854
rect 308048 258586 308368 258618
rect 304674 233778 304706 234334
rect 305262 233778 305294 234334
rect 304674 198334 305294 233778
rect 312114 241774 312734 277218
rect 312114 241218 312146 241774
rect 312702 241218 312734 241774
rect 308048 223174 308368 223206
rect 308048 222938 308090 223174
rect 308326 222938 308368 223174
rect 308048 222854 308368 222938
rect 308048 222618 308090 222854
rect 308326 222618 308368 222854
rect 308048 222586 308368 222618
rect 304674 197778 304706 198334
rect 305262 197778 305294 198334
rect 304674 162334 305294 197778
rect 312114 205774 312734 241218
rect 312114 205218 312146 205774
rect 312702 205218 312734 205774
rect 308048 187174 308368 187206
rect 308048 186938 308090 187174
rect 308326 186938 308368 187174
rect 308048 186854 308368 186938
rect 308048 186618 308090 186854
rect 308326 186618 308368 186854
rect 308048 186586 308368 186618
rect 304674 161778 304706 162334
rect 305262 161778 305294 162334
rect 304674 126334 305294 161778
rect 312114 169774 312734 205218
rect 312114 169218 312146 169774
rect 312702 169218 312734 169774
rect 308048 151174 308368 151206
rect 308048 150938 308090 151174
rect 308326 150938 308368 151174
rect 308048 150854 308368 150938
rect 308048 150618 308090 150854
rect 308326 150618 308368 150854
rect 308048 150586 308368 150618
rect 304674 125778 304706 126334
rect 305262 125778 305294 126334
rect 304674 90334 305294 125778
rect 312114 133774 312734 169218
rect 312114 133218 312146 133774
rect 312702 133218 312734 133774
rect 308048 115174 308368 115206
rect 308048 114938 308090 115174
rect 308326 114938 308368 115174
rect 308048 114854 308368 114938
rect 308048 114618 308090 114854
rect 308326 114618 308368 114854
rect 308048 114586 308368 114618
rect 304674 89778 304706 90334
rect 305262 89778 305294 90334
rect 304674 54334 305294 89778
rect 312114 97774 312734 133218
rect 312114 97218 312146 97774
rect 312702 97218 312734 97774
rect 308048 79174 308368 79206
rect 308048 78938 308090 79174
rect 308326 78938 308368 79174
rect 308048 78854 308368 78938
rect 308048 78618 308090 78854
rect 308326 78618 308368 78854
rect 308048 78586 308368 78618
rect 304674 53778 304706 54334
rect 305262 53778 305294 54334
rect 304674 18334 305294 53778
rect 312114 61774 312734 97218
rect 312114 61218 312146 61774
rect 312702 61218 312734 61774
rect 308048 43174 308368 43206
rect 308048 42938 308090 43174
rect 308326 42938 308368 43174
rect 308048 42854 308368 42938
rect 308048 42618 308090 42854
rect 308326 42618 308368 42854
rect 308048 42586 308368 42618
rect 304674 17778 304706 18334
rect 305262 17778 305294 18334
rect 304674 -4186 305294 17778
rect 312114 25774 312734 61218
rect 312114 25218 312146 25774
rect 312702 25218 312734 25774
rect 308048 7174 308368 7206
rect 308048 6938 308090 7174
rect 308326 6938 308368 7174
rect 308048 6854 308368 6938
rect 308048 6618 308090 6854
rect 308326 6618 308368 6854
rect 308048 6586 308368 6618
rect 304674 -4742 304706 -4186
rect 305262 -4742 305294 -4186
rect 304674 -7654 305294 -4742
rect 312114 -6106 312734 25218
rect 312114 -6662 312146 -6106
rect 312702 -6662 312734 -6106
rect 312114 -7654 312734 -6662
rect 315834 711558 316454 711590
rect 315834 711002 315866 711558
rect 316422 711002 316454 711558
rect 315834 677494 316454 711002
rect 315834 676938 315866 677494
rect 316422 676938 316454 677494
rect 315834 641494 316454 676938
rect 315834 640938 315866 641494
rect 316422 640938 316454 641494
rect 315834 605494 316454 640938
rect 315834 604938 315866 605494
rect 316422 604938 316454 605494
rect 315834 569494 316454 604938
rect 315834 568938 315866 569494
rect 316422 568938 316454 569494
rect 315834 533494 316454 568938
rect 315834 532938 315866 533494
rect 316422 532938 316454 533494
rect 315834 497494 316454 532938
rect 315834 496938 315866 497494
rect 316422 496938 316454 497494
rect 315834 461494 316454 496938
rect 315834 460938 315866 461494
rect 316422 460938 316454 461494
rect 315834 425494 316454 460938
rect 315834 424938 315866 425494
rect 316422 424938 316454 425494
rect 315834 389494 316454 424938
rect 315834 388938 315866 389494
rect 316422 388938 316454 389494
rect 315834 353494 316454 388938
rect 315834 352938 315866 353494
rect 316422 352938 316454 353494
rect 315834 317494 316454 352938
rect 325794 704838 326414 711590
rect 325794 704282 325826 704838
rect 326382 704282 326414 704838
rect 325794 687454 326414 704282
rect 325794 686898 325826 687454
rect 326382 686898 326414 687454
rect 325794 651454 326414 686898
rect 325794 650898 325826 651454
rect 326382 650898 326414 651454
rect 325794 615454 326414 650898
rect 325794 614898 325826 615454
rect 326382 614898 326414 615454
rect 325794 579454 326414 614898
rect 325794 578898 325826 579454
rect 326382 578898 326414 579454
rect 325794 543454 326414 578898
rect 325794 542898 325826 543454
rect 326382 542898 326414 543454
rect 325794 507454 326414 542898
rect 325794 506898 325826 507454
rect 326382 506898 326414 507454
rect 325794 471454 326414 506898
rect 325794 470898 325826 471454
rect 326382 470898 326414 471454
rect 325794 435454 326414 470898
rect 325794 434898 325826 435454
rect 326382 434898 326414 435454
rect 325794 399454 326414 434898
rect 325794 398898 325826 399454
rect 326382 398898 326414 399454
rect 325794 363454 326414 398898
rect 325794 362898 325826 363454
rect 326382 362898 326414 363454
rect 323408 327454 323728 327486
rect 323408 327218 323450 327454
rect 323686 327218 323728 327454
rect 323408 327134 323728 327218
rect 323408 326898 323450 327134
rect 323686 326898 323728 327134
rect 323408 326866 323728 326898
rect 325794 327454 326414 362898
rect 325794 326898 325826 327454
rect 326382 326898 326414 327454
rect 315834 316938 315866 317494
rect 316422 316938 316454 317494
rect 315834 281494 316454 316938
rect 323408 291454 323728 291486
rect 323408 291218 323450 291454
rect 323686 291218 323728 291454
rect 323408 291134 323728 291218
rect 323408 290898 323450 291134
rect 323686 290898 323728 291134
rect 323408 290866 323728 290898
rect 325794 291454 326414 326898
rect 325794 290898 325826 291454
rect 326382 290898 326414 291454
rect 315834 280938 315866 281494
rect 316422 280938 316454 281494
rect 315834 245494 316454 280938
rect 323408 255454 323728 255486
rect 323408 255218 323450 255454
rect 323686 255218 323728 255454
rect 323408 255134 323728 255218
rect 323408 254898 323450 255134
rect 323686 254898 323728 255134
rect 323408 254866 323728 254898
rect 325794 255454 326414 290898
rect 325794 254898 325826 255454
rect 326382 254898 326414 255454
rect 315834 244938 315866 245494
rect 316422 244938 316454 245494
rect 315834 209494 316454 244938
rect 323408 219454 323728 219486
rect 323408 219218 323450 219454
rect 323686 219218 323728 219454
rect 323408 219134 323728 219218
rect 323408 218898 323450 219134
rect 323686 218898 323728 219134
rect 323408 218866 323728 218898
rect 325794 219454 326414 254898
rect 325794 218898 325826 219454
rect 326382 218898 326414 219454
rect 315834 208938 315866 209494
rect 316422 208938 316454 209494
rect 315834 173494 316454 208938
rect 323408 183454 323728 183486
rect 323408 183218 323450 183454
rect 323686 183218 323728 183454
rect 323408 183134 323728 183218
rect 323408 182898 323450 183134
rect 323686 182898 323728 183134
rect 323408 182866 323728 182898
rect 325794 183454 326414 218898
rect 325794 182898 325826 183454
rect 326382 182898 326414 183454
rect 315834 172938 315866 173494
rect 316422 172938 316454 173494
rect 315834 137494 316454 172938
rect 323408 147454 323728 147486
rect 323408 147218 323450 147454
rect 323686 147218 323728 147454
rect 323408 147134 323728 147218
rect 323408 146898 323450 147134
rect 323686 146898 323728 147134
rect 323408 146866 323728 146898
rect 325794 147454 326414 182898
rect 325794 146898 325826 147454
rect 326382 146898 326414 147454
rect 315834 136938 315866 137494
rect 316422 136938 316454 137494
rect 315834 101494 316454 136938
rect 323408 111454 323728 111486
rect 323408 111218 323450 111454
rect 323686 111218 323728 111454
rect 323408 111134 323728 111218
rect 323408 110898 323450 111134
rect 323686 110898 323728 111134
rect 323408 110866 323728 110898
rect 325794 111454 326414 146898
rect 325794 110898 325826 111454
rect 326382 110898 326414 111454
rect 315834 100938 315866 101494
rect 316422 100938 316454 101494
rect 315834 65494 316454 100938
rect 323408 75454 323728 75486
rect 323408 75218 323450 75454
rect 323686 75218 323728 75454
rect 323408 75134 323728 75218
rect 323408 74898 323450 75134
rect 323686 74898 323728 75134
rect 323408 74866 323728 74898
rect 325794 75454 326414 110898
rect 325794 74898 325826 75454
rect 326382 74898 326414 75454
rect 315834 64938 315866 65494
rect 316422 64938 316454 65494
rect 315834 29494 316454 64938
rect 323408 39454 323728 39486
rect 323408 39218 323450 39454
rect 323686 39218 323728 39454
rect 323408 39134 323728 39218
rect 323408 38898 323450 39134
rect 323686 38898 323728 39134
rect 323408 38866 323728 38898
rect 325794 39454 326414 74898
rect 325794 38898 325826 39454
rect 326382 38898 326414 39454
rect 315834 28938 315866 29494
rect 316422 28938 316454 29494
rect 315834 -7066 316454 28938
rect 315834 -7622 315866 -7066
rect 316422 -7622 316454 -7066
rect 315834 -7654 316454 -7622
rect 325794 3454 326414 38898
rect 325794 2898 325826 3454
rect 326382 2898 326414 3454
rect 325794 -346 326414 2898
rect 325794 -902 325826 -346
rect 326382 -902 326414 -346
rect 325794 -7654 326414 -902
rect 329514 705798 330134 711590
rect 329514 705242 329546 705798
rect 330102 705242 330134 705798
rect 329514 691174 330134 705242
rect 329514 690618 329546 691174
rect 330102 690618 330134 691174
rect 329514 655174 330134 690618
rect 329514 654618 329546 655174
rect 330102 654618 330134 655174
rect 329514 619174 330134 654618
rect 329514 618618 329546 619174
rect 330102 618618 330134 619174
rect 329514 583174 330134 618618
rect 329514 582618 329546 583174
rect 330102 582618 330134 583174
rect 329514 547174 330134 582618
rect 329514 546618 329546 547174
rect 330102 546618 330134 547174
rect 329514 511174 330134 546618
rect 329514 510618 329546 511174
rect 330102 510618 330134 511174
rect 329514 475174 330134 510618
rect 329514 474618 329546 475174
rect 330102 474618 330134 475174
rect 329514 439174 330134 474618
rect 329514 438618 329546 439174
rect 330102 438618 330134 439174
rect 329514 403174 330134 438618
rect 329514 402618 329546 403174
rect 330102 402618 330134 403174
rect 329514 367174 330134 402618
rect 329514 366618 329546 367174
rect 330102 366618 330134 367174
rect 329514 331174 330134 366618
rect 329514 330618 329546 331174
rect 330102 330618 330134 331174
rect 329514 295174 330134 330618
rect 329514 294618 329546 295174
rect 330102 294618 330134 295174
rect 329514 259174 330134 294618
rect 329514 258618 329546 259174
rect 330102 258618 330134 259174
rect 329514 223174 330134 258618
rect 329514 222618 329546 223174
rect 330102 222618 330134 223174
rect 329514 187174 330134 222618
rect 329514 186618 329546 187174
rect 330102 186618 330134 187174
rect 329514 151174 330134 186618
rect 329514 150618 329546 151174
rect 330102 150618 330134 151174
rect 329514 115174 330134 150618
rect 329514 114618 329546 115174
rect 330102 114618 330134 115174
rect 329514 79174 330134 114618
rect 329514 78618 329546 79174
rect 330102 78618 330134 79174
rect 329514 43174 330134 78618
rect 329514 42618 329546 43174
rect 330102 42618 330134 43174
rect 329514 7174 330134 42618
rect 329514 6618 329546 7174
rect 330102 6618 330134 7174
rect 329514 -1306 330134 6618
rect 329514 -1862 329546 -1306
rect 330102 -1862 330134 -1306
rect 329514 -7654 330134 -1862
rect 333234 706758 333854 711590
rect 333234 706202 333266 706758
rect 333822 706202 333854 706758
rect 333234 694894 333854 706202
rect 333234 694338 333266 694894
rect 333822 694338 333854 694894
rect 333234 658894 333854 694338
rect 333234 658338 333266 658894
rect 333822 658338 333854 658894
rect 333234 622894 333854 658338
rect 333234 622338 333266 622894
rect 333822 622338 333854 622894
rect 333234 586894 333854 622338
rect 333234 586338 333266 586894
rect 333822 586338 333854 586894
rect 333234 550894 333854 586338
rect 333234 550338 333266 550894
rect 333822 550338 333854 550894
rect 333234 514894 333854 550338
rect 333234 514338 333266 514894
rect 333822 514338 333854 514894
rect 333234 478894 333854 514338
rect 333234 478338 333266 478894
rect 333822 478338 333854 478894
rect 333234 442894 333854 478338
rect 333234 442338 333266 442894
rect 333822 442338 333854 442894
rect 333234 406894 333854 442338
rect 333234 406338 333266 406894
rect 333822 406338 333854 406894
rect 333234 370894 333854 406338
rect 333234 370338 333266 370894
rect 333822 370338 333854 370894
rect 333234 334894 333854 370338
rect 333234 334338 333266 334894
rect 333822 334338 333854 334894
rect 333234 298894 333854 334338
rect 333234 298338 333266 298894
rect 333822 298338 333854 298894
rect 333234 262894 333854 298338
rect 333234 262338 333266 262894
rect 333822 262338 333854 262894
rect 333234 226894 333854 262338
rect 333234 226338 333266 226894
rect 333822 226338 333854 226894
rect 333234 190894 333854 226338
rect 333234 190338 333266 190894
rect 333822 190338 333854 190894
rect 333234 154894 333854 190338
rect 333234 154338 333266 154894
rect 333822 154338 333854 154894
rect 333234 118894 333854 154338
rect 333234 118338 333266 118894
rect 333822 118338 333854 118894
rect 333234 82894 333854 118338
rect 333234 82338 333266 82894
rect 333822 82338 333854 82894
rect 333234 46894 333854 82338
rect 333234 46338 333266 46894
rect 333822 46338 333854 46894
rect 333234 10894 333854 46338
rect 333234 10338 333266 10894
rect 333822 10338 333854 10894
rect 333234 -2266 333854 10338
rect 333234 -2822 333266 -2266
rect 333822 -2822 333854 -2266
rect 333234 -7654 333854 -2822
rect 336954 707718 337574 711590
rect 336954 707162 336986 707718
rect 337542 707162 337574 707718
rect 336954 698614 337574 707162
rect 336954 698058 336986 698614
rect 337542 698058 337574 698614
rect 336954 662614 337574 698058
rect 336954 662058 336986 662614
rect 337542 662058 337574 662614
rect 336954 626614 337574 662058
rect 336954 626058 336986 626614
rect 337542 626058 337574 626614
rect 336954 590614 337574 626058
rect 336954 590058 336986 590614
rect 337542 590058 337574 590614
rect 336954 554614 337574 590058
rect 336954 554058 336986 554614
rect 337542 554058 337574 554614
rect 336954 518614 337574 554058
rect 336954 518058 336986 518614
rect 337542 518058 337574 518614
rect 336954 482614 337574 518058
rect 336954 482058 336986 482614
rect 337542 482058 337574 482614
rect 336954 446614 337574 482058
rect 336954 446058 336986 446614
rect 337542 446058 337574 446614
rect 336954 410614 337574 446058
rect 336954 410058 336986 410614
rect 337542 410058 337574 410614
rect 336954 374614 337574 410058
rect 336954 374058 336986 374614
rect 337542 374058 337574 374614
rect 336954 338614 337574 374058
rect 336954 338058 336986 338614
rect 337542 338058 337574 338614
rect 336954 302614 337574 338058
rect 340674 708678 341294 711590
rect 340674 708122 340706 708678
rect 341262 708122 341294 708678
rect 340674 666334 341294 708122
rect 340674 665778 340706 666334
rect 341262 665778 341294 666334
rect 340674 630334 341294 665778
rect 340674 629778 340706 630334
rect 341262 629778 341294 630334
rect 340674 594334 341294 629778
rect 340674 593778 340706 594334
rect 341262 593778 341294 594334
rect 340674 558334 341294 593778
rect 340674 557778 340706 558334
rect 341262 557778 341294 558334
rect 340674 522334 341294 557778
rect 340674 521778 340706 522334
rect 341262 521778 341294 522334
rect 340674 486334 341294 521778
rect 340674 485778 340706 486334
rect 341262 485778 341294 486334
rect 340674 450334 341294 485778
rect 340674 449778 340706 450334
rect 341262 449778 341294 450334
rect 340674 414334 341294 449778
rect 340674 413778 340706 414334
rect 341262 413778 341294 414334
rect 340674 378334 341294 413778
rect 340674 377778 340706 378334
rect 341262 377778 341294 378334
rect 340674 342334 341294 377778
rect 340674 341778 340706 342334
rect 341262 341778 341294 342334
rect 338768 331174 339088 331206
rect 338768 330938 338810 331174
rect 339046 330938 339088 331174
rect 338768 330854 339088 330938
rect 338768 330618 338810 330854
rect 339046 330618 339088 330854
rect 338768 330586 339088 330618
rect 336954 302058 336986 302614
rect 337542 302058 337574 302614
rect 336954 266614 337574 302058
rect 340674 306334 341294 341778
rect 340674 305778 340706 306334
rect 341262 305778 341294 306334
rect 338768 295174 339088 295206
rect 338768 294938 338810 295174
rect 339046 294938 339088 295174
rect 338768 294854 339088 294938
rect 338768 294618 338810 294854
rect 339046 294618 339088 294854
rect 338768 294586 339088 294618
rect 336954 266058 336986 266614
rect 337542 266058 337574 266614
rect 336954 230614 337574 266058
rect 340674 270334 341294 305778
rect 340674 269778 340706 270334
rect 341262 269778 341294 270334
rect 338768 259174 339088 259206
rect 338768 258938 338810 259174
rect 339046 258938 339088 259174
rect 338768 258854 339088 258938
rect 338768 258618 338810 258854
rect 339046 258618 339088 258854
rect 338768 258586 339088 258618
rect 336954 230058 336986 230614
rect 337542 230058 337574 230614
rect 336954 194614 337574 230058
rect 340674 234334 341294 269778
rect 340674 233778 340706 234334
rect 341262 233778 341294 234334
rect 338768 223174 339088 223206
rect 338768 222938 338810 223174
rect 339046 222938 339088 223174
rect 338768 222854 339088 222938
rect 338768 222618 338810 222854
rect 339046 222618 339088 222854
rect 338768 222586 339088 222618
rect 336954 194058 336986 194614
rect 337542 194058 337574 194614
rect 336954 158614 337574 194058
rect 340674 198334 341294 233778
rect 340674 197778 340706 198334
rect 341262 197778 341294 198334
rect 338768 187174 339088 187206
rect 338768 186938 338810 187174
rect 339046 186938 339088 187174
rect 338768 186854 339088 186938
rect 338768 186618 338810 186854
rect 339046 186618 339088 186854
rect 338768 186586 339088 186618
rect 336954 158058 336986 158614
rect 337542 158058 337574 158614
rect 336954 122614 337574 158058
rect 340674 162334 341294 197778
rect 340674 161778 340706 162334
rect 341262 161778 341294 162334
rect 338768 151174 339088 151206
rect 338768 150938 338810 151174
rect 339046 150938 339088 151174
rect 338768 150854 339088 150938
rect 338768 150618 338810 150854
rect 339046 150618 339088 150854
rect 338768 150586 339088 150618
rect 336954 122058 336986 122614
rect 337542 122058 337574 122614
rect 336954 86614 337574 122058
rect 340674 126334 341294 161778
rect 340674 125778 340706 126334
rect 341262 125778 341294 126334
rect 338768 115174 339088 115206
rect 338768 114938 338810 115174
rect 339046 114938 339088 115174
rect 338768 114854 339088 114938
rect 338768 114618 338810 114854
rect 339046 114618 339088 114854
rect 338768 114586 339088 114618
rect 336954 86058 336986 86614
rect 337542 86058 337574 86614
rect 336954 50614 337574 86058
rect 340674 90334 341294 125778
rect 340674 89778 340706 90334
rect 341262 89778 341294 90334
rect 338768 79174 339088 79206
rect 338768 78938 338810 79174
rect 339046 78938 339088 79174
rect 338768 78854 339088 78938
rect 338768 78618 338810 78854
rect 339046 78618 339088 78854
rect 338768 78586 339088 78618
rect 336954 50058 336986 50614
rect 337542 50058 337574 50614
rect 336954 14614 337574 50058
rect 340674 54334 341294 89778
rect 340674 53778 340706 54334
rect 341262 53778 341294 54334
rect 338768 43174 339088 43206
rect 338768 42938 338810 43174
rect 339046 42938 339088 43174
rect 338768 42854 339088 42938
rect 338768 42618 338810 42854
rect 339046 42618 339088 42854
rect 338768 42586 339088 42618
rect 336954 14058 336986 14614
rect 337542 14058 337574 14614
rect 336954 -3226 337574 14058
rect 340674 18334 341294 53778
rect 340674 17778 340706 18334
rect 341262 17778 341294 18334
rect 338768 7174 339088 7206
rect 338768 6938 338810 7174
rect 339046 6938 339088 7174
rect 338768 6854 339088 6938
rect 338768 6618 338810 6854
rect 339046 6618 339088 6854
rect 338768 6586 339088 6618
rect 336954 -3782 336986 -3226
rect 337542 -3782 337574 -3226
rect 336954 -7654 337574 -3782
rect 340674 -4186 341294 17778
rect 340674 -4742 340706 -4186
rect 341262 -4742 341294 -4186
rect 340674 -7654 341294 -4742
rect 344394 709638 345014 711590
rect 344394 709082 344426 709638
rect 344982 709082 345014 709638
rect 344394 670054 345014 709082
rect 344394 669498 344426 670054
rect 344982 669498 345014 670054
rect 344394 634054 345014 669498
rect 344394 633498 344426 634054
rect 344982 633498 345014 634054
rect 344394 598054 345014 633498
rect 344394 597498 344426 598054
rect 344982 597498 345014 598054
rect 344394 562054 345014 597498
rect 344394 561498 344426 562054
rect 344982 561498 345014 562054
rect 344394 526054 345014 561498
rect 344394 525498 344426 526054
rect 344982 525498 345014 526054
rect 344394 490054 345014 525498
rect 344394 489498 344426 490054
rect 344982 489498 345014 490054
rect 344394 454054 345014 489498
rect 344394 453498 344426 454054
rect 344982 453498 345014 454054
rect 344394 418054 345014 453498
rect 344394 417498 344426 418054
rect 344982 417498 345014 418054
rect 344394 382054 345014 417498
rect 344394 381498 344426 382054
rect 344982 381498 345014 382054
rect 344394 346054 345014 381498
rect 344394 345498 344426 346054
rect 344982 345498 345014 346054
rect 344394 310054 345014 345498
rect 344394 309498 344426 310054
rect 344982 309498 345014 310054
rect 344394 274054 345014 309498
rect 344394 273498 344426 274054
rect 344982 273498 345014 274054
rect 344394 238054 345014 273498
rect 344394 237498 344426 238054
rect 344982 237498 345014 238054
rect 344394 202054 345014 237498
rect 344394 201498 344426 202054
rect 344982 201498 345014 202054
rect 344394 166054 345014 201498
rect 344394 165498 344426 166054
rect 344982 165498 345014 166054
rect 344394 130054 345014 165498
rect 344394 129498 344426 130054
rect 344982 129498 345014 130054
rect 344394 94054 345014 129498
rect 344394 93498 344426 94054
rect 344982 93498 345014 94054
rect 344394 58054 345014 93498
rect 344394 57498 344426 58054
rect 344982 57498 345014 58054
rect 344394 22054 345014 57498
rect 344394 21498 344426 22054
rect 344982 21498 345014 22054
rect 344394 -5146 345014 21498
rect 344394 -5702 344426 -5146
rect 344982 -5702 345014 -5146
rect 344394 -7654 345014 -5702
rect 348114 710598 348734 711590
rect 348114 710042 348146 710598
rect 348702 710042 348734 710598
rect 348114 673774 348734 710042
rect 348114 673218 348146 673774
rect 348702 673218 348734 673774
rect 348114 637774 348734 673218
rect 348114 637218 348146 637774
rect 348702 637218 348734 637774
rect 348114 601774 348734 637218
rect 348114 601218 348146 601774
rect 348702 601218 348734 601774
rect 348114 565774 348734 601218
rect 348114 565218 348146 565774
rect 348702 565218 348734 565774
rect 348114 529774 348734 565218
rect 348114 529218 348146 529774
rect 348702 529218 348734 529774
rect 348114 493774 348734 529218
rect 348114 493218 348146 493774
rect 348702 493218 348734 493774
rect 348114 457774 348734 493218
rect 348114 457218 348146 457774
rect 348702 457218 348734 457774
rect 348114 421774 348734 457218
rect 348114 421218 348146 421774
rect 348702 421218 348734 421774
rect 348114 385774 348734 421218
rect 348114 385218 348146 385774
rect 348702 385218 348734 385774
rect 348114 349774 348734 385218
rect 348114 349218 348146 349774
rect 348702 349218 348734 349774
rect 348114 313774 348734 349218
rect 348114 313218 348146 313774
rect 348702 313218 348734 313774
rect 348114 277774 348734 313218
rect 348114 277218 348146 277774
rect 348702 277218 348734 277774
rect 348114 241774 348734 277218
rect 348114 241218 348146 241774
rect 348702 241218 348734 241774
rect 348114 205774 348734 241218
rect 348114 205218 348146 205774
rect 348702 205218 348734 205774
rect 348114 169774 348734 205218
rect 348114 169218 348146 169774
rect 348702 169218 348734 169774
rect 348114 133774 348734 169218
rect 348114 133218 348146 133774
rect 348702 133218 348734 133774
rect 348114 97774 348734 133218
rect 348114 97218 348146 97774
rect 348702 97218 348734 97774
rect 348114 61774 348734 97218
rect 348114 61218 348146 61774
rect 348702 61218 348734 61774
rect 348114 25774 348734 61218
rect 348114 25218 348146 25774
rect 348702 25218 348734 25774
rect 348114 -6106 348734 25218
rect 348114 -6662 348146 -6106
rect 348702 -6662 348734 -6106
rect 348114 -7654 348734 -6662
rect 351834 711558 352454 711590
rect 351834 711002 351866 711558
rect 352422 711002 352454 711558
rect 351834 677494 352454 711002
rect 351834 676938 351866 677494
rect 352422 676938 352454 677494
rect 351834 641494 352454 676938
rect 351834 640938 351866 641494
rect 352422 640938 352454 641494
rect 351834 605494 352454 640938
rect 351834 604938 351866 605494
rect 352422 604938 352454 605494
rect 351834 569494 352454 604938
rect 351834 568938 351866 569494
rect 352422 568938 352454 569494
rect 351834 533494 352454 568938
rect 351834 532938 351866 533494
rect 352422 532938 352454 533494
rect 351834 497494 352454 532938
rect 351834 496938 351866 497494
rect 352422 496938 352454 497494
rect 351834 461494 352454 496938
rect 351834 460938 351866 461494
rect 352422 460938 352454 461494
rect 351834 425494 352454 460938
rect 351834 424938 351866 425494
rect 352422 424938 352454 425494
rect 351834 389494 352454 424938
rect 351834 388938 351866 389494
rect 352422 388938 352454 389494
rect 351834 353494 352454 388938
rect 351834 352938 351866 353494
rect 352422 352938 352454 353494
rect 351834 317494 352454 352938
rect 361794 704838 362414 711590
rect 361794 704282 361826 704838
rect 362382 704282 362414 704838
rect 361794 687454 362414 704282
rect 361794 686898 361826 687454
rect 362382 686898 362414 687454
rect 361794 651454 362414 686898
rect 361794 650898 361826 651454
rect 362382 650898 362414 651454
rect 361794 615454 362414 650898
rect 361794 614898 361826 615454
rect 362382 614898 362414 615454
rect 361794 579454 362414 614898
rect 361794 578898 361826 579454
rect 362382 578898 362414 579454
rect 361794 543454 362414 578898
rect 361794 542898 361826 543454
rect 362382 542898 362414 543454
rect 361794 507454 362414 542898
rect 361794 506898 361826 507454
rect 362382 506898 362414 507454
rect 361794 471454 362414 506898
rect 361794 470898 361826 471454
rect 362382 470898 362414 471454
rect 361794 435454 362414 470898
rect 361794 434898 361826 435454
rect 362382 434898 362414 435454
rect 361794 399454 362414 434898
rect 361794 398898 361826 399454
rect 362382 398898 362414 399454
rect 361794 363454 362414 398898
rect 361794 362898 361826 363454
rect 362382 362898 362414 363454
rect 354128 327454 354448 327486
rect 354128 327218 354170 327454
rect 354406 327218 354448 327454
rect 354128 327134 354448 327218
rect 354128 326898 354170 327134
rect 354406 326898 354448 327134
rect 354128 326866 354448 326898
rect 361794 327454 362414 362898
rect 361794 326898 361826 327454
rect 362382 326898 362414 327454
rect 351834 316938 351866 317494
rect 352422 316938 352454 317494
rect 351834 281494 352454 316938
rect 354128 291454 354448 291486
rect 354128 291218 354170 291454
rect 354406 291218 354448 291454
rect 354128 291134 354448 291218
rect 354128 290898 354170 291134
rect 354406 290898 354448 291134
rect 354128 290866 354448 290898
rect 361794 291454 362414 326898
rect 361794 290898 361826 291454
rect 362382 290898 362414 291454
rect 351834 280938 351866 281494
rect 352422 280938 352454 281494
rect 351834 245494 352454 280938
rect 354128 255454 354448 255486
rect 354128 255218 354170 255454
rect 354406 255218 354448 255454
rect 354128 255134 354448 255218
rect 354128 254898 354170 255134
rect 354406 254898 354448 255134
rect 354128 254866 354448 254898
rect 361794 255454 362414 290898
rect 361794 254898 361826 255454
rect 362382 254898 362414 255454
rect 351834 244938 351866 245494
rect 352422 244938 352454 245494
rect 351834 209494 352454 244938
rect 354128 219454 354448 219486
rect 354128 219218 354170 219454
rect 354406 219218 354448 219454
rect 354128 219134 354448 219218
rect 354128 218898 354170 219134
rect 354406 218898 354448 219134
rect 354128 218866 354448 218898
rect 361794 219454 362414 254898
rect 361794 218898 361826 219454
rect 362382 218898 362414 219454
rect 351834 208938 351866 209494
rect 352422 208938 352454 209494
rect 351834 173494 352454 208938
rect 354128 183454 354448 183486
rect 354128 183218 354170 183454
rect 354406 183218 354448 183454
rect 354128 183134 354448 183218
rect 354128 182898 354170 183134
rect 354406 182898 354448 183134
rect 354128 182866 354448 182898
rect 361794 183454 362414 218898
rect 361794 182898 361826 183454
rect 362382 182898 362414 183454
rect 351834 172938 351866 173494
rect 352422 172938 352454 173494
rect 351834 137494 352454 172938
rect 354128 147454 354448 147486
rect 354128 147218 354170 147454
rect 354406 147218 354448 147454
rect 354128 147134 354448 147218
rect 354128 146898 354170 147134
rect 354406 146898 354448 147134
rect 354128 146866 354448 146898
rect 361794 147454 362414 182898
rect 361794 146898 361826 147454
rect 362382 146898 362414 147454
rect 351834 136938 351866 137494
rect 352422 136938 352454 137494
rect 351834 101494 352454 136938
rect 354128 111454 354448 111486
rect 354128 111218 354170 111454
rect 354406 111218 354448 111454
rect 354128 111134 354448 111218
rect 354128 110898 354170 111134
rect 354406 110898 354448 111134
rect 354128 110866 354448 110898
rect 361794 111454 362414 146898
rect 361794 110898 361826 111454
rect 362382 110898 362414 111454
rect 351834 100938 351866 101494
rect 352422 100938 352454 101494
rect 351834 65494 352454 100938
rect 354128 75454 354448 75486
rect 354128 75218 354170 75454
rect 354406 75218 354448 75454
rect 354128 75134 354448 75218
rect 354128 74898 354170 75134
rect 354406 74898 354448 75134
rect 354128 74866 354448 74898
rect 361794 75454 362414 110898
rect 361794 74898 361826 75454
rect 362382 74898 362414 75454
rect 351834 64938 351866 65494
rect 352422 64938 352454 65494
rect 351834 29494 352454 64938
rect 354128 39454 354448 39486
rect 354128 39218 354170 39454
rect 354406 39218 354448 39454
rect 354128 39134 354448 39218
rect 354128 38898 354170 39134
rect 354406 38898 354448 39134
rect 354128 38866 354448 38898
rect 361794 39454 362414 74898
rect 361794 38898 361826 39454
rect 362382 38898 362414 39454
rect 351834 28938 351866 29494
rect 352422 28938 352454 29494
rect 351834 -7066 352454 28938
rect 351834 -7622 351866 -7066
rect 352422 -7622 352454 -7066
rect 351834 -7654 352454 -7622
rect 361794 3454 362414 38898
rect 361794 2898 361826 3454
rect 362382 2898 362414 3454
rect 365514 705798 366134 711590
rect 365514 705242 365546 705798
rect 366102 705242 366134 705798
rect 365514 691174 366134 705242
rect 365514 690618 365546 691174
rect 366102 690618 366134 691174
rect 365514 655174 366134 690618
rect 365514 654618 365546 655174
rect 366102 654618 366134 655174
rect 365514 619174 366134 654618
rect 365514 618618 365546 619174
rect 366102 618618 366134 619174
rect 365514 583174 366134 618618
rect 365514 582618 365546 583174
rect 366102 582618 366134 583174
rect 365514 547174 366134 582618
rect 365514 546618 365546 547174
rect 366102 546618 366134 547174
rect 365514 511174 366134 546618
rect 365514 510618 365546 511174
rect 366102 510618 366134 511174
rect 365514 475174 366134 510618
rect 365514 474618 365546 475174
rect 366102 474618 366134 475174
rect 365514 439174 366134 474618
rect 365514 438618 365546 439174
rect 366102 438618 366134 439174
rect 365514 403174 366134 438618
rect 365514 402618 365546 403174
rect 366102 402618 366134 403174
rect 365514 367174 366134 402618
rect 365514 366618 365546 367174
rect 366102 366618 366134 367174
rect 365514 331174 366134 366618
rect 369234 706758 369854 711590
rect 369234 706202 369266 706758
rect 369822 706202 369854 706758
rect 369234 694894 369854 706202
rect 369234 694338 369266 694894
rect 369822 694338 369854 694894
rect 369234 658894 369854 694338
rect 369234 658338 369266 658894
rect 369822 658338 369854 658894
rect 369234 622894 369854 658338
rect 369234 622338 369266 622894
rect 369822 622338 369854 622894
rect 369234 586894 369854 622338
rect 369234 586338 369266 586894
rect 369822 586338 369854 586894
rect 369234 550894 369854 586338
rect 369234 550338 369266 550894
rect 369822 550338 369854 550894
rect 369234 514894 369854 550338
rect 369234 514338 369266 514894
rect 369822 514338 369854 514894
rect 369234 478894 369854 514338
rect 369234 478338 369266 478894
rect 369822 478338 369854 478894
rect 369234 442894 369854 478338
rect 369234 442338 369266 442894
rect 369822 442338 369854 442894
rect 369234 406894 369854 442338
rect 369234 406338 369266 406894
rect 369822 406338 369854 406894
rect 369234 370894 369854 406338
rect 369234 370338 369266 370894
rect 369822 370338 369854 370894
rect 369234 354980 369854 370338
rect 372954 707718 373574 711590
rect 372954 707162 372986 707718
rect 373542 707162 373574 707718
rect 372954 698614 373574 707162
rect 372954 698058 372986 698614
rect 373542 698058 373574 698614
rect 372954 662614 373574 698058
rect 372954 662058 372986 662614
rect 373542 662058 373574 662614
rect 372954 626614 373574 662058
rect 372954 626058 372986 626614
rect 373542 626058 373574 626614
rect 372954 590614 373574 626058
rect 372954 590058 372986 590614
rect 373542 590058 373574 590614
rect 372954 554614 373574 590058
rect 372954 554058 372986 554614
rect 373542 554058 373574 554614
rect 372954 518614 373574 554058
rect 372954 518058 372986 518614
rect 373542 518058 373574 518614
rect 372954 482614 373574 518058
rect 372954 482058 372986 482614
rect 373542 482058 373574 482614
rect 372954 446614 373574 482058
rect 372954 446058 372986 446614
rect 373542 446058 373574 446614
rect 372954 410614 373574 446058
rect 372954 410058 372986 410614
rect 373542 410058 373574 410614
rect 372954 374614 373574 410058
rect 372954 374058 372986 374614
rect 373542 374058 373574 374614
rect 372954 338614 373574 374058
rect 372954 338058 372986 338614
rect 373542 338058 373574 338614
rect 365514 330618 365546 331174
rect 366102 330618 366134 331174
rect 365514 295174 366134 330618
rect 369488 331174 369808 331206
rect 369488 330938 369530 331174
rect 369766 330938 369808 331174
rect 369488 330854 369808 330938
rect 369488 330618 369530 330854
rect 369766 330618 369808 330854
rect 369488 330586 369808 330618
rect 372954 302614 373574 338058
rect 372954 302058 372986 302614
rect 373542 302058 373574 302614
rect 365514 294618 365546 295174
rect 366102 294618 366134 295174
rect 365514 259174 366134 294618
rect 369488 295174 369808 295206
rect 369488 294938 369530 295174
rect 369766 294938 369808 295174
rect 369488 294854 369808 294938
rect 369488 294618 369530 294854
rect 369766 294618 369808 294854
rect 369488 294586 369808 294618
rect 372954 266614 373574 302058
rect 372954 266058 372986 266614
rect 373542 266058 373574 266614
rect 365514 258618 365546 259174
rect 366102 258618 366134 259174
rect 365514 223174 366134 258618
rect 369488 259174 369808 259206
rect 369488 258938 369530 259174
rect 369766 258938 369808 259174
rect 369488 258854 369808 258938
rect 369488 258618 369530 258854
rect 369766 258618 369808 258854
rect 369488 258586 369808 258618
rect 372954 230614 373574 266058
rect 372954 230058 372986 230614
rect 373542 230058 373574 230614
rect 365514 222618 365546 223174
rect 366102 222618 366134 223174
rect 365514 187174 366134 222618
rect 369488 223174 369808 223206
rect 369488 222938 369530 223174
rect 369766 222938 369808 223174
rect 369488 222854 369808 222938
rect 369488 222618 369530 222854
rect 369766 222618 369808 222854
rect 369488 222586 369808 222618
rect 372954 194614 373574 230058
rect 372954 194058 372986 194614
rect 373542 194058 373574 194614
rect 365514 186618 365546 187174
rect 366102 186618 366134 187174
rect 365514 151174 366134 186618
rect 369488 187174 369808 187206
rect 369488 186938 369530 187174
rect 369766 186938 369808 187174
rect 369488 186854 369808 186938
rect 369488 186618 369530 186854
rect 369766 186618 369808 186854
rect 369488 186586 369808 186618
rect 372954 158614 373574 194058
rect 372954 158058 372986 158614
rect 373542 158058 373574 158614
rect 365514 150618 365546 151174
rect 366102 150618 366134 151174
rect 365514 115174 366134 150618
rect 369488 151174 369808 151206
rect 369488 150938 369530 151174
rect 369766 150938 369808 151174
rect 369488 150854 369808 150938
rect 369488 150618 369530 150854
rect 369766 150618 369808 150854
rect 369488 150586 369808 150618
rect 372954 122614 373574 158058
rect 372954 122058 372986 122614
rect 373542 122058 373574 122614
rect 365514 114618 365546 115174
rect 366102 114618 366134 115174
rect 365514 79174 366134 114618
rect 369488 115174 369808 115206
rect 369488 114938 369530 115174
rect 369766 114938 369808 115174
rect 369488 114854 369808 114938
rect 369488 114618 369530 114854
rect 369766 114618 369808 114854
rect 369488 114586 369808 114618
rect 372954 86614 373574 122058
rect 372954 86058 372986 86614
rect 373542 86058 373574 86614
rect 365514 78618 365546 79174
rect 366102 78618 366134 79174
rect 365514 43174 366134 78618
rect 369488 79174 369808 79206
rect 369488 78938 369530 79174
rect 369766 78938 369808 79174
rect 369488 78854 369808 78938
rect 369488 78618 369530 78854
rect 369766 78618 369808 78854
rect 369488 78586 369808 78618
rect 372954 50614 373574 86058
rect 372954 50058 372986 50614
rect 373542 50058 373574 50614
rect 365514 42618 365546 43174
rect 366102 42618 366134 43174
rect 365514 7174 366134 42618
rect 369488 43174 369808 43206
rect 369488 42938 369530 43174
rect 369766 42938 369808 43174
rect 369488 42854 369808 42938
rect 369488 42618 369530 42854
rect 369766 42618 369808 42854
rect 369488 42586 369808 42618
rect 372954 14614 373574 50058
rect 372954 14058 372986 14614
rect 373542 14058 373574 14614
rect 365514 6618 365546 7174
rect 366102 6618 366134 7174
rect 364195 3092 364261 3093
rect 364195 3028 364196 3092
rect 364260 3028 364261 3092
rect 364195 3027 364261 3028
rect 361794 -346 362414 2898
rect 364198 2821 364258 3027
rect 364195 2820 364261 2821
rect 364195 2756 364196 2820
rect 364260 2756 364261 2820
rect 364195 2755 364261 2756
rect 361794 -902 361826 -346
rect 362382 -902 362414 -346
rect 361794 -7654 362414 -902
rect 365514 -1306 366134 6618
rect 369488 7174 369808 7206
rect 369488 6938 369530 7174
rect 369766 6938 369808 7174
rect 369488 6854 369808 6938
rect 369488 6618 369530 6854
rect 369766 6618 369808 6854
rect 369488 6586 369808 6618
rect 365514 -1862 365546 -1306
rect 366102 -1862 366134 -1306
rect 365514 -7654 366134 -1862
rect 372954 -3226 373574 14058
rect 372954 -3782 372986 -3226
rect 373542 -3782 373574 -3226
rect 372954 -7654 373574 -3782
rect 376674 708678 377294 711590
rect 376674 708122 376706 708678
rect 377262 708122 377294 708678
rect 376674 666334 377294 708122
rect 376674 665778 376706 666334
rect 377262 665778 377294 666334
rect 376674 630334 377294 665778
rect 376674 629778 376706 630334
rect 377262 629778 377294 630334
rect 376674 594334 377294 629778
rect 376674 593778 376706 594334
rect 377262 593778 377294 594334
rect 376674 558334 377294 593778
rect 376674 557778 376706 558334
rect 377262 557778 377294 558334
rect 376674 522334 377294 557778
rect 376674 521778 376706 522334
rect 377262 521778 377294 522334
rect 376674 486334 377294 521778
rect 376674 485778 376706 486334
rect 377262 485778 377294 486334
rect 376674 450334 377294 485778
rect 376674 449778 376706 450334
rect 377262 449778 377294 450334
rect 376674 414334 377294 449778
rect 376674 413778 376706 414334
rect 377262 413778 377294 414334
rect 376674 378334 377294 413778
rect 376674 377778 376706 378334
rect 377262 377778 377294 378334
rect 376674 342334 377294 377778
rect 376674 341778 376706 342334
rect 377262 341778 377294 342334
rect 376674 306334 377294 341778
rect 376674 305778 376706 306334
rect 377262 305778 377294 306334
rect 376674 270334 377294 305778
rect 376674 269778 376706 270334
rect 377262 269778 377294 270334
rect 376674 234334 377294 269778
rect 376674 233778 376706 234334
rect 377262 233778 377294 234334
rect 376674 198334 377294 233778
rect 376674 197778 376706 198334
rect 377262 197778 377294 198334
rect 376674 162334 377294 197778
rect 376674 161778 376706 162334
rect 377262 161778 377294 162334
rect 376674 126334 377294 161778
rect 376674 125778 376706 126334
rect 377262 125778 377294 126334
rect 376674 90334 377294 125778
rect 376674 89778 376706 90334
rect 377262 89778 377294 90334
rect 376674 54334 377294 89778
rect 376674 53778 376706 54334
rect 377262 53778 377294 54334
rect 376674 18334 377294 53778
rect 376674 17778 376706 18334
rect 377262 17778 377294 18334
rect 376674 -4186 377294 17778
rect 380394 709638 381014 711590
rect 380394 709082 380426 709638
rect 380982 709082 381014 709638
rect 380394 670054 381014 709082
rect 380394 669498 380426 670054
rect 380982 669498 381014 670054
rect 380394 634054 381014 669498
rect 380394 633498 380426 634054
rect 380982 633498 381014 634054
rect 380394 598054 381014 633498
rect 380394 597498 380426 598054
rect 380982 597498 381014 598054
rect 380394 562054 381014 597498
rect 380394 561498 380426 562054
rect 380982 561498 381014 562054
rect 380394 526054 381014 561498
rect 380394 525498 380426 526054
rect 380982 525498 381014 526054
rect 380394 490054 381014 525498
rect 380394 489498 380426 490054
rect 380982 489498 381014 490054
rect 380394 454054 381014 489498
rect 380394 453498 380426 454054
rect 380982 453498 381014 454054
rect 380394 418054 381014 453498
rect 380394 417498 380426 418054
rect 380982 417498 381014 418054
rect 380394 382054 381014 417498
rect 380394 381498 380426 382054
rect 380982 381498 381014 382054
rect 380394 346054 381014 381498
rect 384114 710598 384734 711590
rect 384114 710042 384146 710598
rect 384702 710042 384734 710598
rect 384114 673774 384734 710042
rect 384114 673218 384146 673774
rect 384702 673218 384734 673774
rect 384114 637774 384734 673218
rect 384114 637218 384146 637774
rect 384702 637218 384734 637774
rect 384114 601774 384734 637218
rect 384114 601218 384146 601774
rect 384702 601218 384734 601774
rect 384114 565774 384734 601218
rect 384114 565218 384146 565774
rect 384702 565218 384734 565774
rect 384114 529774 384734 565218
rect 384114 529218 384146 529774
rect 384702 529218 384734 529774
rect 384114 493774 384734 529218
rect 384114 493218 384146 493774
rect 384702 493218 384734 493774
rect 384114 457774 384734 493218
rect 384114 457218 384146 457774
rect 384702 457218 384734 457774
rect 384114 421774 384734 457218
rect 384114 421218 384146 421774
rect 384702 421218 384734 421774
rect 384114 385774 384734 421218
rect 384114 385218 384146 385774
rect 384702 385218 384734 385774
rect 384114 354980 384734 385218
rect 387834 711558 388454 711590
rect 387834 711002 387866 711558
rect 388422 711002 388454 711558
rect 387834 677494 388454 711002
rect 387834 676938 387866 677494
rect 388422 676938 388454 677494
rect 387834 641494 388454 676938
rect 387834 640938 387866 641494
rect 388422 640938 388454 641494
rect 387834 605494 388454 640938
rect 387834 604938 387866 605494
rect 388422 604938 388454 605494
rect 387834 569494 388454 604938
rect 387834 568938 387866 569494
rect 388422 568938 388454 569494
rect 387834 533494 388454 568938
rect 387834 532938 387866 533494
rect 388422 532938 388454 533494
rect 387834 497494 388454 532938
rect 387834 496938 387866 497494
rect 388422 496938 388454 497494
rect 387834 461494 388454 496938
rect 387834 460938 387866 461494
rect 388422 460938 388454 461494
rect 387834 425494 388454 460938
rect 387834 424938 387866 425494
rect 388422 424938 388454 425494
rect 387834 389494 388454 424938
rect 387834 388938 387866 389494
rect 388422 388938 388454 389494
rect 380394 345498 380426 346054
rect 380982 345498 381014 346054
rect 380394 310054 381014 345498
rect 387834 353494 388454 388938
rect 387834 352938 387866 353494
rect 388422 352938 388454 353494
rect 384848 327454 385168 327486
rect 384848 327218 384890 327454
rect 385126 327218 385168 327454
rect 384848 327134 385168 327218
rect 384848 326898 384890 327134
rect 385126 326898 385168 327134
rect 384848 326866 385168 326898
rect 380394 309498 380426 310054
rect 380982 309498 381014 310054
rect 380394 274054 381014 309498
rect 387834 317494 388454 352938
rect 387834 316938 387866 317494
rect 388422 316938 388454 317494
rect 384848 291454 385168 291486
rect 384848 291218 384890 291454
rect 385126 291218 385168 291454
rect 384848 291134 385168 291218
rect 384848 290898 384890 291134
rect 385126 290898 385168 291134
rect 384848 290866 385168 290898
rect 380394 273498 380426 274054
rect 380982 273498 381014 274054
rect 380394 238054 381014 273498
rect 387834 281494 388454 316938
rect 387834 280938 387866 281494
rect 388422 280938 388454 281494
rect 384848 255454 385168 255486
rect 384848 255218 384890 255454
rect 385126 255218 385168 255454
rect 384848 255134 385168 255218
rect 384848 254898 384890 255134
rect 385126 254898 385168 255134
rect 384848 254866 385168 254898
rect 380394 237498 380426 238054
rect 380982 237498 381014 238054
rect 380394 202054 381014 237498
rect 387834 245494 388454 280938
rect 387834 244938 387866 245494
rect 388422 244938 388454 245494
rect 384848 219454 385168 219486
rect 384848 219218 384890 219454
rect 385126 219218 385168 219454
rect 384848 219134 385168 219218
rect 384848 218898 384890 219134
rect 385126 218898 385168 219134
rect 384848 218866 385168 218898
rect 380394 201498 380426 202054
rect 380982 201498 381014 202054
rect 380394 166054 381014 201498
rect 387834 209494 388454 244938
rect 387834 208938 387866 209494
rect 388422 208938 388454 209494
rect 384848 183454 385168 183486
rect 384848 183218 384890 183454
rect 385126 183218 385168 183454
rect 384848 183134 385168 183218
rect 384848 182898 384890 183134
rect 385126 182898 385168 183134
rect 384848 182866 385168 182898
rect 380394 165498 380426 166054
rect 380982 165498 381014 166054
rect 380394 130054 381014 165498
rect 387834 173494 388454 208938
rect 387834 172938 387866 173494
rect 388422 172938 388454 173494
rect 384848 147454 385168 147486
rect 384848 147218 384890 147454
rect 385126 147218 385168 147454
rect 384848 147134 385168 147218
rect 384848 146898 384890 147134
rect 385126 146898 385168 147134
rect 384848 146866 385168 146898
rect 380394 129498 380426 130054
rect 380982 129498 381014 130054
rect 380394 94054 381014 129498
rect 387834 137494 388454 172938
rect 387834 136938 387866 137494
rect 388422 136938 388454 137494
rect 384848 111454 385168 111486
rect 384848 111218 384890 111454
rect 385126 111218 385168 111454
rect 384848 111134 385168 111218
rect 384848 110898 384890 111134
rect 385126 110898 385168 111134
rect 384848 110866 385168 110898
rect 380394 93498 380426 94054
rect 380982 93498 381014 94054
rect 380394 58054 381014 93498
rect 387834 101494 388454 136938
rect 387834 100938 387866 101494
rect 388422 100938 388454 101494
rect 384848 75454 385168 75486
rect 384848 75218 384890 75454
rect 385126 75218 385168 75454
rect 384848 75134 385168 75218
rect 384848 74898 384890 75134
rect 385126 74898 385168 75134
rect 384848 74866 385168 74898
rect 380394 57498 380426 58054
rect 380982 57498 381014 58054
rect 380394 22054 381014 57498
rect 387834 65494 388454 100938
rect 387834 64938 387866 65494
rect 388422 64938 388454 65494
rect 384848 39454 385168 39486
rect 384848 39218 384890 39454
rect 385126 39218 385168 39454
rect 384848 39134 385168 39218
rect 384848 38898 384890 39134
rect 385126 38898 385168 39134
rect 384848 38866 385168 38898
rect 380394 21498 380426 22054
rect 380982 21498 381014 22054
rect 377443 3092 377509 3093
rect 377443 3028 377444 3092
rect 377508 3028 377509 3092
rect 377443 3027 377509 3028
rect 377446 2549 377506 3027
rect 377443 2548 377509 2549
rect 377443 2484 377444 2548
rect 377508 2484 377509 2548
rect 377443 2483 377509 2484
rect 376674 -4742 376706 -4186
rect 377262 -4742 377294 -4186
rect 376674 -7654 377294 -4742
rect 380394 -5146 381014 21498
rect 387834 29494 388454 64938
rect 387834 28938 387866 29494
rect 388422 28938 388454 29494
rect 383515 3772 383581 3773
rect 383515 3708 383516 3772
rect 383580 3708 383581 3772
rect 383515 3707 383581 3708
rect 383518 2549 383578 3707
rect 383515 2548 383581 2549
rect 383515 2484 383516 2548
rect 383580 2484 383581 2548
rect 383515 2483 383581 2484
rect 380394 -5702 380426 -5146
rect 380982 -5702 381014 -5146
rect 380394 -7654 381014 -5702
rect 387834 -7066 388454 28938
rect 397794 704838 398414 711590
rect 397794 704282 397826 704838
rect 398382 704282 398414 704838
rect 397794 687454 398414 704282
rect 397794 686898 397826 687454
rect 398382 686898 398414 687454
rect 397794 651454 398414 686898
rect 397794 650898 397826 651454
rect 398382 650898 398414 651454
rect 397794 615454 398414 650898
rect 397794 614898 397826 615454
rect 398382 614898 398414 615454
rect 397794 579454 398414 614898
rect 397794 578898 397826 579454
rect 398382 578898 398414 579454
rect 397794 543454 398414 578898
rect 397794 542898 397826 543454
rect 398382 542898 398414 543454
rect 397794 507454 398414 542898
rect 397794 506898 397826 507454
rect 398382 506898 398414 507454
rect 397794 471454 398414 506898
rect 397794 470898 397826 471454
rect 398382 470898 398414 471454
rect 397794 435454 398414 470898
rect 397794 434898 397826 435454
rect 398382 434898 398414 435454
rect 397794 399454 398414 434898
rect 397794 398898 397826 399454
rect 398382 398898 398414 399454
rect 397794 363454 398414 398898
rect 397794 362898 397826 363454
rect 398382 362898 398414 363454
rect 397794 327454 398414 362898
rect 401514 705798 402134 711590
rect 401514 705242 401546 705798
rect 402102 705242 402134 705798
rect 401514 691174 402134 705242
rect 401514 690618 401546 691174
rect 402102 690618 402134 691174
rect 401514 655174 402134 690618
rect 401514 654618 401546 655174
rect 402102 654618 402134 655174
rect 401514 619174 402134 654618
rect 401514 618618 401546 619174
rect 402102 618618 402134 619174
rect 401514 583174 402134 618618
rect 401514 582618 401546 583174
rect 402102 582618 402134 583174
rect 401514 547174 402134 582618
rect 401514 546618 401546 547174
rect 402102 546618 402134 547174
rect 401514 511174 402134 546618
rect 401514 510618 401546 511174
rect 402102 510618 402134 511174
rect 401514 475174 402134 510618
rect 401514 474618 401546 475174
rect 402102 474618 402134 475174
rect 401514 439174 402134 474618
rect 401514 438618 401546 439174
rect 402102 438618 402134 439174
rect 401514 403174 402134 438618
rect 401514 402618 401546 403174
rect 402102 402618 402134 403174
rect 401514 367174 402134 402618
rect 401514 366618 401546 367174
rect 402102 366618 402134 367174
rect 400208 331174 400528 331206
rect 400208 330938 400250 331174
rect 400486 330938 400528 331174
rect 400208 330854 400528 330938
rect 400208 330618 400250 330854
rect 400486 330618 400528 330854
rect 400208 330586 400528 330618
rect 401514 331174 402134 366618
rect 401514 330618 401546 331174
rect 402102 330618 402134 331174
rect 397794 326898 397826 327454
rect 398382 326898 398414 327454
rect 397794 291454 398414 326898
rect 400208 295174 400528 295206
rect 400208 294938 400250 295174
rect 400486 294938 400528 295174
rect 400208 294854 400528 294938
rect 400208 294618 400250 294854
rect 400486 294618 400528 294854
rect 400208 294586 400528 294618
rect 401514 295174 402134 330618
rect 401514 294618 401546 295174
rect 402102 294618 402134 295174
rect 397794 290898 397826 291454
rect 398382 290898 398414 291454
rect 397794 255454 398414 290898
rect 400208 259174 400528 259206
rect 400208 258938 400250 259174
rect 400486 258938 400528 259174
rect 400208 258854 400528 258938
rect 400208 258618 400250 258854
rect 400486 258618 400528 258854
rect 400208 258586 400528 258618
rect 401514 259174 402134 294618
rect 401514 258618 401546 259174
rect 402102 258618 402134 259174
rect 397794 254898 397826 255454
rect 398382 254898 398414 255454
rect 397794 219454 398414 254898
rect 400208 223174 400528 223206
rect 400208 222938 400250 223174
rect 400486 222938 400528 223174
rect 400208 222854 400528 222938
rect 400208 222618 400250 222854
rect 400486 222618 400528 222854
rect 400208 222586 400528 222618
rect 401514 223174 402134 258618
rect 401514 222618 401546 223174
rect 402102 222618 402134 223174
rect 397794 218898 397826 219454
rect 398382 218898 398414 219454
rect 397794 183454 398414 218898
rect 400208 187174 400528 187206
rect 400208 186938 400250 187174
rect 400486 186938 400528 187174
rect 400208 186854 400528 186938
rect 400208 186618 400250 186854
rect 400486 186618 400528 186854
rect 400208 186586 400528 186618
rect 401514 187174 402134 222618
rect 401514 186618 401546 187174
rect 402102 186618 402134 187174
rect 397794 182898 397826 183454
rect 398382 182898 398414 183454
rect 397794 147454 398414 182898
rect 400208 151174 400528 151206
rect 400208 150938 400250 151174
rect 400486 150938 400528 151174
rect 400208 150854 400528 150938
rect 400208 150618 400250 150854
rect 400486 150618 400528 150854
rect 400208 150586 400528 150618
rect 401514 151174 402134 186618
rect 401514 150618 401546 151174
rect 402102 150618 402134 151174
rect 397794 146898 397826 147454
rect 398382 146898 398414 147454
rect 397794 111454 398414 146898
rect 400208 115174 400528 115206
rect 400208 114938 400250 115174
rect 400486 114938 400528 115174
rect 400208 114854 400528 114938
rect 400208 114618 400250 114854
rect 400486 114618 400528 114854
rect 400208 114586 400528 114618
rect 401514 115174 402134 150618
rect 401514 114618 401546 115174
rect 402102 114618 402134 115174
rect 397794 110898 397826 111454
rect 398382 110898 398414 111454
rect 397794 75454 398414 110898
rect 400208 79174 400528 79206
rect 400208 78938 400250 79174
rect 400486 78938 400528 79174
rect 400208 78854 400528 78938
rect 400208 78618 400250 78854
rect 400486 78618 400528 78854
rect 400208 78586 400528 78618
rect 401514 79174 402134 114618
rect 401514 78618 401546 79174
rect 402102 78618 402134 79174
rect 397794 74898 397826 75454
rect 398382 74898 398414 75454
rect 397794 39454 398414 74898
rect 400208 43174 400528 43206
rect 400208 42938 400250 43174
rect 400486 42938 400528 43174
rect 400208 42854 400528 42938
rect 400208 42618 400250 42854
rect 400486 42618 400528 42854
rect 400208 42586 400528 42618
rect 401514 43174 402134 78618
rect 401514 42618 401546 43174
rect 402102 42618 402134 43174
rect 397794 38898 397826 39454
rect 398382 38898 398414 39454
rect 389403 3772 389469 3773
rect 389403 3708 389404 3772
rect 389468 3708 389469 3772
rect 389403 3707 389469 3708
rect 389406 2549 389466 3707
rect 397794 3454 398414 38898
rect 400208 7174 400528 7206
rect 400208 6938 400250 7174
rect 400486 6938 400528 7174
rect 400208 6854 400528 6938
rect 400208 6618 400250 6854
rect 400486 6618 400528 6854
rect 400208 6586 400528 6618
rect 401514 7174 402134 42618
rect 401514 6618 401546 7174
rect 402102 6618 402134 7174
rect 397499 3364 397565 3365
rect 397499 3300 397500 3364
rect 397564 3300 397565 3364
rect 397499 3299 397565 3300
rect 397502 2685 397562 3299
rect 397794 2898 397826 3454
rect 398382 2898 398414 3454
rect 397499 2684 397565 2685
rect 397499 2620 397500 2684
rect 397564 2620 397565 2684
rect 397499 2619 397565 2620
rect 389403 2548 389469 2549
rect 389403 2484 389404 2548
rect 389468 2484 389469 2548
rect 389403 2483 389469 2484
rect 387834 -7622 387866 -7066
rect 388422 -7622 388454 -7066
rect 387834 -7654 388454 -7622
rect 397794 -346 398414 2898
rect 397794 -902 397826 -346
rect 398382 -902 398414 -346
rect 397794 -7654 398414 -902
rect 401514 -1306 402134 6618
rect 401514 -1862 401546 -1306
rect 402102 -1862 402134 -1306
rect 401514 -7654 402134 -1862
rect 405234 706758 405854 711590
rect 405234 706202 405266 706758
rect 405822 706202 405854 706758
rect 405234 694894 405854 706202
rect 405234 694338 405266 694894
rect 405822 694338 405854 694894
rect 405234 658894 405854 694338
rect 405234 658338 405266 658894
rect 405822 658338 405854 658894
rect 405234 622894 405854 658338
rect 405234 622338 405266 622894
rect 405822 622338 405854 622894
rect 405234 586894 405854 622338
rect 405234 586338 405266 586894
rect 405822 586338 405854 586894
rect 405234 550894 405854 586338
rect 405234 550338 405266 550894
rect 405822 550338 405854 550894
rect 405234 514894 405854 550338
rect 405234 514338 405266 514894
rect 405822 514338 405854 514894
rect 405234 478894 405854 514338
rect 405234 478338 405266 478894
rect 405822 478338 405854 478894
rect 405234 442894 405854 478338
rect 405234 442338 405266 442894
rect 405822 442338 405854 442894
rect 405234 406894 405854 442338
rect 405234 406338 405266 406894
rect 405822 406338 405854 406894
rect 405234 370894 405854 406338
rect 405234 370338 405266 370894
rect 405822 370338 405854 370894
rect 405234 334894 405854 370338
rect 405234 334338 405266 334894
rect 405822 334338 405854 334894
rect 405234 298894 405854 334338
rect 405234 298338 405266 298894
rect 405822 298338 405854 298894
rect 405234 262894 405854 298338
rect 405234 262338 405266 262894
rect 405822 262338 405854 262894
rect 405234 226894 405854 262338
rect 405234 226338 405266 226894
rect 405822 226338 405854 226894
rect 405234 190894 405854 226338
rect 405234 190338 405266 190894
rect 405822 190338 405854 190894
rect 405234 154894 405854 190338
rect 405234 154338 405266 154894
rect 405822 154338 405854 154894
rect 405234 118894 405854 154338
rect 405234 118338 405266 118894
rect 405822 118338 405854 118894
rect 405234 82894 405854 118338
rect 405234 82338 405266 82894
rect 405822 82338 405854 82894
rect 405234 46894 405854 82338
rect 405234 46338 405266 46894
rect 405822 46338 405854 46894
rect 405234 10894 405854 46338
rect 405234 10338 405266 10894
rect 405822 10338 405854 10894
rect 405234 -2266 405854 10338
rect 408954 707718 409574 711590
rect 408954 707162 408986 707718
rect 409542 707162 409574 707718
rect 408954 698614 409574 707162
rect 408954 698058 408986 698614
rect 409542 698058 409574 698614
rect 408954 662614 409574 698058
rect 408954 662058 408986 662614
rect 409542 662058 409574 662614
rect 408954 626614 409574 662058
rect 408954 626058 408986 626614
rect 409542 626058 409574 626614
rect 408954 590614 409574 626058
rect 408954 590058 408986 590614
rect 409542 590058 409574 590614
rect 408954 554614 409574 590058
rect 408954 554058 408986 554614
rect 409542 554058 409574 554614
rect 408954 518614 409574 554058
rect 408954 518058 408986 518614
rect 409542 518058 409574 518614
rect 408954 482614 409574 518058
rect 408954 482058 408986 482614
rect 409542 482058 409574 482614
rect 408954 446614 409574 482058
rect 408954 446058 408986 446614
rect 409542 446058 409574 446614
rect 408954 410614 409574 446058
rect 408954 410058 408986 410614
rect 409542 410058 409574 410614
rect 408954 374614 409574 410058
rect 408954 374058 408986 374614
rect 409542 374058 409574 374614
rect 408954 338614 409574 374058
rect 408954 338058 408986 338614
rect 409542 338058 409574 338614
rect 408954 302614 409574 338058
rect 408954 302058 408986 302614
rect 409542 302058 409574 302614
rect 408954 266614 409574 302058
rect 408954 266058 408986 266614
rect 409542 266058 409574 266614
rect 408954 230614 409574 266058
rect 408954 230058 408986 230614
rect 409542 230058 409574 230614
rect 408954 194614 409574 230058
rect 408954 194058 408986 194614
rect 409542 194058 409574 194614
rect 408954 158614 409574 194058
rect 408954 158058 408986 158614
rect 409542 158058 409574 158614
rect 408954 122614 409574 158058
rect 408954 122058 408986 122614
rect 409542 122058 409574 122614
rect 408954 86614 409574 122058
rect 408954 86058 408986 86614
rect 409542 86058 409574 86614
rect 408954 50614 409574 86058
rect 408954 50058 408986 50614
rect 409542 50058 409574 50614
rect 408954 14614 409574 50058
rect 408954 14058 408986 14614
rect 409542 14058 409574 14614
rect 405963 3228 406029 3229
rect 405963 3164 405964 3228
rect 406028 3164 406029 3228
rect 405963 3163 406029 3164
rect 405966 2821 406026 3163
rect 405963 2820 406029 2821
rect 405963 2756 405964 2820
rect 406028 2756 406029 2820
rect 405963 2755 406029 2756
rect 405234 -2822 405266 -2266
rect 405822 -2822 405854 -2266
rect 405234 -7654 405854 -2822
rect 408954 -3226 409574 14058
rect 408954 -3782 408986 -3226
rect 409542 -3782 409574 -3226
rect 408954 -7654 409574 -3782
rect 412674 708678 413294 711590
rect 412674 708122 412706 708678
rect 413262 708122 413294 708678
rect 412674 666334 413294 708122
rect 412674 665778 412706 666334
rect 413262 665778 413294 666334
rect 412674 630334 413294 665778
rect 412674 629778 412706 630334
rect 413262 629778 413294 630334
rect 412674 594334 413294 629778
rect 412674 593778 412706 594334
rect 413262 593778 413294 594334
rect 412674 558334 413294 593778
rect 412674 557778 412706 558334
rect 413262 557778 413294 558334
rect 412674 522334 413294 557778
rect 412674 521778 412706 522334
rect 413262 521778 413294 522334
rect 412674 486334 413294 521778
rect 412674 485778 412706 486334
rect 413262 485778 413294 486334
rect 412674 450334 413294 485778
rect 412674 449778 412706 450334
rect 413262 449778 413294 450334
rect 412674 414334 413294 449778
rect 412674 413778 412706 414334
rect 413262 413778 413294 414334
rect 412674 378334 413294 413778
rect 412674 377778 412706 378334
rect 413262 377778 413294 378334
rect 412674 342334 413294 377778
rect 412674 341778 412706 342334
rect 413262 341778 413294 342334
rect 412674 306334 413294 341778
rect 416394 709638 417014 711590
rect 416394 709082 416426 709638
rect 416982 709082 417014 709638
rect 416394 670054 417014 709082
rect 416394 669498 416426 670054
rect 416982 669498 417014 670054
rect 416394 634054 417014 669498
rect 416394 633498 416426 634054
rect 416982 633498 417014 634054
rect 416394 598054 417014 633498
rect 416394 597498 416426 598054
rect 416982 597498 417014 598054
rect 416394 562054 417014 597498
rect 416394 561498 416426 562054
rect 416982 561498 417014 562054
rect 416394 526054 417014 561498
rect 416394 525498 416426 526054
rect 416982 525498 417014 526054
rect 416394 490054 417014 525498
rect 416394 489498 416426 490054
rect 416982 489498 417014 490054
rect 416394 454054 417014 489498
rect 416394 453498 416426 454054
rect 416982 453498 417014 454054
rect 416394 418054 417014 453498
rect 416394 417498 416426 418054
rect 416982 417498 417014 418054
rect 416394 382054 417014 417498
rect 416394 381498 416426 382054
rect 416982 381498 417014 382054
rect 416394 346054 417014 381498
rect 416394 345498 416426 346054
rect 416982 345498 417014 346054
rect 415568 327454 415888 327486
rect 415568 327218 415610 327454
rect 415846 327218 415888 327454
rect 415568 327134 415888 327218
rect 415568 326898 415610 327134
rect 415846 326898 415888 327134
rect 415568 326866 415888 326898
rect 412674 305778 412706 306334
rect 413262 305778 413294 306334
rect 412674 270334 413294 305778
rect 416394 310054 417014 345498
rect 416394 309498 416426 310054
rect 416982 309498 417014 310054
rect 415568 291454 415888 291486
rect 415568 291218 415610 291454
rect 415846 291218 415888 291454
rect 415568 291134 415888 291218
rect 415568 290898 415610 291134
rect 415846 290898 415888 291134
rect 415568 290866 415888 290898
rect 412674 269778 412706 270334
rect 413262 269778 413294 270334
rect 412674 234334 413294 269778
rect 416394 274054 417014 309498
rect 416394 273498 416426 274054
rect 416982 273498 417014 274054
rect 415568 255454 415888 255486
rect 415568 255218 415610 255454
rect 415846 255218 415888 255454
rect 415568 255134 415888 255218
rect 415568 254898 415610 255134
rect 415846 254898 415888 255134
rect 415568 254866 415888 254898
rect 412674 233778 412706 234334
rect 413262 233778 413294 234334
rect 412674 198334 413294 233778
rect 416394 238054 417014 273498
rect 416394 237498 416426 238054
rect 416982 237498 417014 238054
rect 415568 219454 415888 219486
rect 415568 219218 415610 219454
rect 415846 219218 415888 219454
rect 415568 219134 415888 219218
rect 415568 218898 415610 219134
rect 415846 218898 415888 219134
rect 415568 218866 415888 218898
rect 412674 197778 412706 198334
rect 413262 197778 413294 198334
rect 412674 162334 413294 197778
rect 416394 202054 417014 237498
rect 416394 201498 416426 202054
rect 416982 201498 417014 202054
rect 415568 183454 415888 183486
rect 415568 183218 415610 183454
rect 415846 183218 415888 183454
rect 415568 183134 415888 183218
rect 415568 182898 415610 183134
rect 415846 182898 415888 183134
rect 415568 182866 415888 182898
rect 412674 161778 412706 162334
rect 413262 161778 413294 162334
rect 412674 126334 413294 161778
rect 416394 166054 417014 201498
rect 416394 165498 416426 166054
rect 416982 165498 417014 166054
rect 415568 147454 415888 147486
rect 415568 147218 415610 147454
rect 415846 147218 415888 147454
rect 415568 147134 415888 147218
rect 415568 146898 415610 147134
rect 415846 146898 415888 147134
rect 415568 146866 415888 146898
rect 412674 125778 412706 126334
rect 413262 125778 413294 126334
rect 412674 90334 413294 125778
rect 416394 130054 417014 165498
rect 416394 129498 416426 130054
rect 416982 129498 417014 130054
rect 415568 111454 415888 111486
rect 415568 111218 415610 111454
rect 415846 111218 415888 111454
rect 415568 111134 415888 111218
rect 415568 110898 415610 111134
rect 415846 110898 415888 111134
rect 415568 110866 415888 110898
rect 412674 89778 412706 90334
rect 413262 89778 413294 90334
rect 412674 54334 413294 89778
rect 416394 94054 417014 129498
rect 416394 93498 416426 94054
rect 416982 93498 417014 94054
rect 415568 75454 415888 75486
rect 415568 75218 415610 75454
rect 415846 75218 415888 75454
rect 415568 75134 415888 75218
rect 415568 74898 415610 75134
rect 415846 74898 415888 75134
rect 415568 74866 415888 74898
rect 412674 53778 412706 54334
rect 413262 53778 413294 54334
rect 412674 18334 413294 53778
rect 416394 58054 417014 93498
rect 416394 57498 416426 58054
rect 416982 57498 417014 58054
rect 415568 39454 415888 39486
rect 415568 39218 415610 39454
rect 415846 39218 415888 39454
rect 415568 39134 415888 39218
rect 415568 38898 415610 39134
rect 415846 38898 415888 39134
rect 415568 38866 415888 38898
rect 412674 17778 412706 18334
rect 413262 17778 413294 18334
rect 412674 -4186 413294 17778
rect 412674 -4742 412706 -4186
rect 413262 -4742 413294 -4186
rect 412674 -7654 413294 -4742
rect 416394 22054 417014 57498
rect 416394 21498 416426 22054
rect 416982 21498 417014 22054
rect 416394 -5146 417014 21498
rect 416394 -5702 416426 -5146
rect 416982 -5702 417014 -5146
rect 416394 -7654 417014 -5702
rect 420114 710598 420734 711590
rect 420114 710042 420146 710598
rect 420702 710042 420734 710598
rect 420114 673774 420734 710042
rect 420114 673218 420146 673774
rect 420702 673218 420734 673774
rect 420114 637774 420734 673218
rect 420114 637218 420146 637774
rect 420702 637218 420734 637774
rect 420114 601774 420734 637218
rect 420114 601218 420146 601774
rect 420702 601218 420734 601774
rect 420114 565774 420734 601218
rect 420114 565218 420146 565774
rect 420702 565218 420734 565774
rect 420114 529774 420734 565218
rect 420114 529218 420146 529774
rect 420702 529218 420734 529774
rect 420114 493774 420734 529218
rect 420114 493218 420146 493774
rect 420702 493218 420734 493774
rect 420114 457774 420734 493218
rect 420114 457218 420146 457774
rect 420702 457218 420734 457774
rect 420114 421774 420734 457218
rect 420114 421218 420146 421774
rect 420702 421218 420734 421774
rect 420114 385774 420734 421218
rect 420114 385218 420146 385774
rect 420702 385218 420734 385774
rect 420114 349774 420734 385218
rect 420114 349218 420146 349774
rect 420702 349218 420734 349774
rect 420114 313774 420734 349218
rect 420114 313218 420146 313774
rect 420702 313218 420734 313774
rect 420114 277774 420734 313218
rect 420114 277218 420146 277774
rect 420702 277218 420734 277774
rect 420114 241774 420734 277218
rect 420114 241218 420146 241774
rect 420702 241218 420734 241774
rect 420114 205774 420734 241218
rect 420114 205218 420146 205774
rect 420702 205218 420734 205774
rect 420114 169774 420734 205218
rect 420114 169218 420146 169774
rect 420702 169218 420734 169774
rect 420114 133774 420734 169218
rect 420114 133218 420146 133774
rect 420702 133218 420734 133774
rect 420114 97774 420734 133218
rect 420114 97218 420146 97774
rect 420702 97218 420734 97774
rect 420114 61774 420734 97218
rect 420114 61218 420146 61774
rect 420702 61218 420734 61774
rect 420114 25774 420734 61218
rect 420114 25218 420146 25774
rect 420702 25218 420734 25774
rect 420114 -6106 420734 25218
rect 420114 -6662 420146 -6106
rect 420702 -6662 420734 -6106
rect 420114 -7654 420734 -6662
rect 423834 711558 424454 711590
rect 423834 711002 423866 711558
rect 424422 711002 424454 711558
rect 423834 677494 424454 711002
rect 423834 676938 423866 677494
rect 424422 676938 424454 677494
rect 423834 641494 424454 676938
rect 423834 640938 423866 641494
rect 424422 640938 424454 641494
rect 423834 605494 424454 640938
rect 423834 604938 423866 605494
rect 424422 604938 424454 605494
rect 423834 569494 424454 604938
rect 423834 568938 423866 569494
rect 424422 568938 424454 569494
rect 423834 533494 424454 568938
rect 423834 532938 423866 533494
rect 424422 532938 424454 533494
rect 423834 497494 424454 532938
rect 423834 496938 423866 497494
rect 424422 496938 424454 497494
rect 423834 461494 424454 496938
rect 423834 460938 423866 461494
rect 424422 460938 424454 461494
rect 423834 425494 424454 460938
rect 423834 424938 423866 425494
rect 424422 424938 424454 425494
rect 423834 389494 424454 424938
rect 423834 388938 423866 389494
rect 424422 388938 424454 389494
rect 423834 353494 424454 388938
rect 423834 352938 423866 353494
rect 424422 352938 424454 353494
rect 423834 317494 424454 352938
rect 433794 704838 434414 711590
rect 433794 704282 433826 704838
rect 434382 704282 434414 704838
rect 433794 687454 434414 704282
rect 433794 686898 433826 687454
rect 434382 686898 434414 687454
rect 433794 651454 434414 686898
rect 433794 650898 433826 651454
rect 434382 650898 434414 651454
rect 433794 615454 434414 650898
rect 433794 614898 433826 615454
rect 434382 614898 434414 615454
rect 433794 579454 434414 614898
rect 433794 578898 433826 579454
rect 434382 578898 434414 579454
rect 433794 543454 434414 578898
rect 433794 542898 433826 543454
rect 434382 542898 434414 543454
rect 433794 507454 434414 542898
rect 433794 506898 433826 507454
rect 434382 506898 434414 507454
rect 433794 471454 434414 506898
rect 433794 470898 433826 471454
rect 434382 470898 434414 471454
rect 433794 435454 434414 470898
rect 433794 434898 433826 435454
rect 434382 434898 434414 435454
rect 433794 399454 434414 434898
rect 433794 398898 433826 399454
rect 434382 398898 434414 399454
rect 433794 363454 434414 398898
rect 433794 362898 433826 363454
rect 434382 362898 434414 363454
rect 430928 331174 431248 331206
rect 430928 330938 430970 331174
rect 431206 330938 431248 331174
rect 430928 330854 431248 330938
rect 430928 330618 430970 330854
rect 431206 330618 431248 330854
rect 430928 330586 431248 330618
rect 423834 316938 423866 317494
rect 424422 316938 424454 317494
rect 423834 281494 424454 316938
rect 433794 327454 434414 362898
rect 433794 326898 433826 327454
rect 434382 326898 434414 327454
rect 430928 295174 431248 295206
rect 430928 294938 430970 295174
rect 431206 294938 431248 295174
rect 430928 294854 431248 294938
rect 430928 294618 430970 294854
rect 431206 294618 431248 294854
rect 430928 294586 431248 294618
rect 423834 280938 423866 281494
rect 424422 280938 424454 281494
rect 423834 245494 424454 280938
rect 433794 291454 434414 326898
rect 433794 290898 433826 291454
rect 434382 290898 434414 291454
rect 430928 259174 431248 259206
rect 430928 258938 430970 259174
rect 431206 258938 431248 259174
rect 430928 258854 431248 258938
rect 430928 258618 430970 258854
rect 431206 258618 431248 258854
rect 430928 258586 431248 258618
rect 423834 244938 423866 245494
rect 424422 244938 424454 245494
rect 423834 209494 424454 244938
rect 433794 255454 434414 290898
rect 433794 254898 433826 255454
rect 434382 254898 434414 255454
rect 430928 223174 431248 223206
rect 430928 222938 430970 223174
rect 431206 222938 431248 223174
rect 430928 222854 431248 222938
rect 430928 222618 430970 222854
rect 431206 222618 431248 222854
rect 430928 222586 431248 222618
rect 423834 208938 423866 209494
rect 424422 208938 424454 209494
rect 423834 173494 424454 208938
rect 433794 219454 434414 254898
rect 433794 218898 433826 219454
rect 434382 218898 434414 219454
rect 430928 187174 431248 187206
rect 430928 186938 430970 187174
rect 431206 186938 431248 187174
rect 430928 186854 431248 186938
rect 430928 186618 430970 186854
rect 431206 186618 431248 186854
rect 430928 186586 431248 186618
rect 423834 172938 423866 173494
rect 424422 172938 424454 173494
rect 423834 137494 424454 172938
rect 433794 183454 434414 218898
rect 433794 182898 433826 183454
rect 434382 182898 434414 183454
rect 430928 151174 431248 151206
rect 430928 150938 430970 151174
rect 431206 150938 431248 151174
rect 430928 150854 431248 150938
rect 430928 150618 430970 150854
rect 431206 150618 431248 150854
rect 430928 150586 431248 150618
rect 423834 136938 423866 137494
rect 424422 136938 424454 137494
rect 423834 101494 424454 136938
rect 433794 147454 434414 182898
rect 433794 146898 433826 147454
rect 434382 146898 434414 147454
rect 430928 115174 431248 115206
rect 430928 114938 430970 115174
rect 431206 114938 431248 115174
rect 430928 114854 431248 114938
rect 430928 114618 430970 114854
rect 431206 114618 431248 114854
rect 430928 114586 431248 114618
rect 423834 100938 423866 101494
rect 424422 100938 424454 101494
rect 423834 65494 424454 100938
rect 433794 111454 434414 146898
rect 433794 110898 433826 111454
rect 434382 110898 434414 111454
rect 430928 79174 431248 79206
rect 430928 78938 430970 79174
rect 431206 78938 431248 79174
rect 430928 78854 431248 78938
rect 430928 78618 430970 78854
rect 431206 78618 431248 78854
rect 430928 78586 431248 78618
rect 423834 64938 423866 65494
rect 424422 64938 424454 65494
rect 423834 29494 424454 64938
rect 433794 75454 434414 110898
rect 433794 74898 433826 75454
rect 434382 74898 434414 75454
rect 430928 43174 431248 43206
rect 430928 42938 430970 43174
rect 431206 42938 431248 43174
rect 430928 42854 431248 42938
rect 430928 42618 430970 42854
rect 431206 42618 431248 42854
rect 430928 42586 431248 42618
rect 423834 28938 423866 29494
rect 424422 28938 424454 29494
rect 423834 -7066 424454 28938
rect 433794 39454 434414 74898
rect 433794 38898 433826 39454
rect 434382 38898 434414 39454
rect 430928 7174 431248 7206
rect 430928 6938 430970 7174
rect 431206 6938 431248 7174
rect 430928 6854 431248 6938
rect 430928 6618 430970 6854
rect 431206 6618 431248 6854
rect 430928 6586 431248 6618
rect 423834 -7622 423866 -7066
rect 424422 -7622 424454 -7066
rect 423834 -7654 424454 -7622
rect 433794 3454 434414 38898
rect 433794 2898 433826 3454
rect 434382 2898 434414 3454
rect 433794 -346 434414 2898
rect 433794 -902 433826 -346
rect 434382 -902 434414 -346
rect 433794 -7654 434414 -902
rect 437514 705798 438134 711590
rect 437514 705242 437546 705798
rect 438102 705242 438134 705798
rect 437514 691174 438134 705242
rect 437514 690618 437546 691174
rect 438102 690618 438134 691174
rect 437514 655174 438134 690618
rect 437514 654618 437546 655174
rect 438102 654618 438134 655174
rect 437514 619174 438134 654618
rect 437514 618618 437546 619174
rect 438102 618618 438134 619174
rect 437514 583174 438134 618618
rect 437514 582618 437546 583174
rect 438102 582618 438134 583174
rect 437514 547174 438134 582618
rect 437514 546618 437546 547174
rect 438102 546618 438134 547174
rect 437514 511174 438134 546618
rect 437514 510618 437546 511174
rect 438102 510618 438134 511174
rect 437514 475174 438134 510618
rect 437514 474618 437546 475174
rect 438102 474618 438134 475174
rect 437514 439174 438134 474618
rect 437514 438618 437546 439174
rect 438102 438618 438134 439174
rect 437514 403174 438134 438618
rect 437514 402618 437546 403174
rect 438102 402618 438134 403174
rect 437514 367174 438134 402618
rect 437514 366618 437546 367174
rect 438102 366618 438134 367174
rect 437514 331174 438134 366618
rect 437514 330618 437546 331174
rect 438102 330618 438134 331174
rect 437514 295174 438134 330618
rect 437514 294618 437546 295174
rect 438102 294618 438134 295174
rect 437514 259174 438134 294618
rect 437514 258618 437546 259174
rect 438102 258618 438134 259174
rect 437514 223174 438134 258618
rect 437514 222618 437546 223174
rect 438102 222618 438134 223174
rect 437514 187174 438134 222618
rect 437514 186618 437546 187174
rect 438102 186618 438134 187174
rect 437514 151174 438134 186618
rect 437514 150618 437546 151174
rect 438102 150618 438134 151174
rect 437514 115174 438134 150618
rect 437514 114618 437546 115174
rect 438102 114618 438134 115174
rect 437514 79174 438134 114618
rect 437514 78618 437546 79174
rect 438102 78618 438134 79174
rect 437514 43174 438134 78618
rect 437514 42618 437546 43174
rect 438102 42618 438134 43174
rect 437514 7174 438134 42618
rect 437514 6618 437546 7174
rect 438102 6618 438134 7174
rect 437514 -1306 438134 6618
rect 437514 -1862 437546 -1306
rect 438102 -1862 438134 -1306
rect 437514 -7654 438134 -1862
rect 441234 706758 441854 711590
rect 441234 706202 441266 706758
rect 441822 706202 441854 706758
rect 441234 694894 441854 706202
rect 441234 694338 441266 694894
rect 441822 694338 441854 694894
rect 441234 658894 441854 694338
rect 441234 658338 441266 658894
rect 441822 658338 441854 658894
rect 441234 622894 441854 658338
rect 441234 622338 441266 622894
rect 441822 622338 441854 622894
rect 441234 586894 441854 622338
rect 441234 586338 441266 586894
rect 441822 586338 441854 586894
rect 441234 550894 441854 586338
rect 441234 550338 441266 550894
rect 441822 550338 441854 550894
rect 441234 514894 441854 550338
rect 441234 514338 441266 514894
rect 441822 514338 441854 514894
rect 441234 478894 441854 514338
rect 441234 478338 441266 478894
rect 441822 478338 441854 478894
rect 441234 442894 441854 478338
rect 441234 442338 441266 442894
rect 441822 442338 441854 442894
rect 441234 406894 441854 442338
rect 441234 406338 441266 406894
rect 441822 406338 441854 406894
rect 441234 370894 441854 406338
rect 441234 370338 441266 370894
rect 441822 370338 441854 370894
rect 441234 334894 441854 370338
rect 441234 334338 441266 334894
rect 441822 334338 441854 334894
rect 441234 298894 441854 334338
rect 441234 298338 441266 298894
rect 441822 298338 441854 298894
rect 441234 262894 441854 298338
rect 441234 262338 441266 262894
rect 441822 262338 441854 262894
rect 441234 226894 441854 262338
rect 441234 226338 441266 226894
rect 441822 226338 441854 226894
rect 441234 190894 441854 226338
rect 441234 190338 441266 190894
rect 441822 190338 441854 190894
rect 441234 154894 441854 190338
rect 441234 154338 441266 154894
rect 441822 154338 441854 154894
rect 441234 118894 441854 154338
rect 441234 118338 441266 118894
rect 441822 118338 441854 118894
rect 441234 82894 441854 118338
rect 441234 82338 441266 82894
rect 441822 82338 441854 82894
rect 441234 46894 441854 82338
rect 441234 46338 441266 46894
rect 441822 46338 441854 46894
rect 441234 10894 441854 46338
rect 441234 10338 441266 10894
rect 441822 10338 441854 10894
rect 441234 -2266 441854 10338
rect 441234 -2822 441266 -2266
rect 441822 -2822 441854 -2266
rect 441234 -7654 441854 -2822
rect 444954 707718 445574 711590
rect 444954 707162 444986 707718
rect 445542 707162 445574 707718
rect 444954 698614 445574 707162
rect 444954 698058 444986 698614
rect 445542 698058 445574 698614
rect 444954 662614 445574 698058
rect 444954 662058 444986 662614
rect 445542 662058 445574 662614
rect 444954 626614 445574 662058
rect 444954 626058 444986 626614
rect 445542 626058 445574 626614
rect 444954 590614 445574 626058
rect 444954 590058 444986 590614
rect 445542 590058 445574 590614
rect 444954 554614 445574 590058
rect 444954 554058 444986 554614
rect 445542 554058 445574 554614
rect 444954 518614 445574 554058
rect 444954 518058 444986 518614
rect 445542 518058 445574 518614
rect 444954 482614 445574 518058
rect 444954 482058 444986 482614
rect 445542 482058 445574 482614
rect 444954 446614 445574 482058
rect 444954 446058 444986 446614
rect 445542 446058 445574 446614
rect 444954 410614 445574 446058
rect 444954 410058 444986 410614
rect 445542 410058 445574 410614
rect 444954 374614 445574 410058
rect 444954 374058 444986 374614
rect 445542 374058 445574 374614
rect 444954 338614 445574 374058
rect 444954 338058 444986 338614
rect 445542 338058 445574 338614
rect 444954 302614 445574 338058
rect 448674 708678 449294 711590
rect 448674 708122 448706 708678
rect 449262 708122 449294 708678
rect 448674 666334 449294 708122
rect 448674 665778 448706 666334
rect 449262 665778 449294 666334
rect 448674 630334 449294 665778
rect 448674 629778 448706 630334
rect 449262 629778 449294 630334
rect 448674 594334 449294 629778
rect 448674 593778 448706 594334
rect 449262 593778 449294 594334
rect 448674 558334 449294 593778
rect 448674 557778 448706 558334
rect 449262 557778 449294 558334
rect 448674 522334 449294 557778
rect 448674 521778 448706 522334
rect 449262 521778 449294 522334
rect 448674 486334 449294 521778
rect 448674 485778 448706 486334
rect 449262 485778 449294 486334
rect 448674 450334 449294 485778
rect 448674 449778 448706 450334
rect 449262 449778 449294 450334
rect 448674 414334 449294 449778
rect 448674 413778 448706 414334
rect 449262 413778 449294 414334
rect 448674 378334 449294 413778
rect 448674 377778 448706 378334
rect 449262 377778 449294 378334
rect 448674 342334 449294 377778
rect 448674 341778 448706 342334
rect 449262 341778 449294 342334
rect 446288 327454 446608 327486
rect 446288 327218 446330 327454
rect 446566 327218 446608 327454
rect 446288 327134 446608 327218
rect 446288 326898 446330 327134
rect 446566 326898 446608 327134
rect 446288 326866 446608 326898
rect 444954 302058 444986 302614
rect 445542 302058 445574 302614
rect 444954 266614 445574 302058
rect 448674 306334 449294 341778
rect 448674 305778 448706 306334
rect 449262 305778 449294 306334
rect 446288 291454 446608 291486
rect 446288 291218 446330 291454
rect 446566 291218 446608 291454
rect 446288 291134 446608 291218
rect 446288 290898 446330 291134
rect 446566 290898 446608 291134
rect 446288 290866 446608 290898
rect 444954 266058 444986 266614
rect 445542 266058 445574 266614
rect 444954 230614 445574 266058
rect 448674 270334 449294 305778
rect 448674 269778 448706 270334
rect 449262 269778 449294 270334
rect 446288 255454 446608 255486
rect 446288 255218 446330 255454
rect 446566 255218 446608 255454
rect 446288 255134 446608 255218
rect 446288 254898 446330 255134
rect 446566 254898 446608 255134
rect 446288 254866 446608 254898
rect 444954 230058 444986 230614
rect 445542 230058 445574 230614
rect 444954 194614 445574 230058
rect 448674 234334 449294 269778
rect 448674 233778 448706 234334
rect 449262 233778 449294 234334
rect 446288 219454 446608 219486
rect 446288 219218 446330 219454
rect 446566 219218 446608 219454
rect 446288 219134 446608 219218
rect 446288 218898 446330 219134
rect 446566 218898 446608 219134
rect 446288 218866 446608 218898
rect 444954 194058 444986 194614
rect 445542 194058 445574 194614
rect 444954 158614 445574 194058
rect 448674 198334 449294 233778
rect 448674 197778 448706 198334
rect 449262 197778 449294 198334
rect 446288 183454 446608 183486
rect 446288 183218 446330 183454
rect 446566 183218 446608 183454
rect 446288 183134 446608 183218
rect 446288 182898 446330 183134
rect 446566 182898 446608 183134
rect 446288 182866 446608 182898
rect 444954 158058 444986 158614
rect 445542 158058 445574 158614
rect 444954 122614 445574 158058
rect 448674 162334 449294 197778
rect 448674 161778 448706 162334
rect 449262 161778 449294 162334
rect 446288 147454 446608 147486
rect 446288 147218 446330 147454
rect 446566 147218 446608 147454
rect 446288 147134 446608 147218
rect 446288 146898 446330 147134
rect 446566 146898 446608 147134
rect 446288 146866 446608 146898
rect 444954 122058 444986 122614
rect 445542 122058 445574 122614
rect 444954 86614 445574 122058
rect 448674 126334 449294 161778
rect 448674 125778 448706 126334
rect 449262 125778 449294 126334
rect 446288 111454 446608 111486
rect 446288 111218 446330 111454
rect 446566 111218 446608 111454
rect 446288 111134 446608 111218
rect 446288 110898 446330 111134
rect 446566 110898 446608 111134
rect 446288 110866 446608 110898
rect 444954 86058 444986 86614
rect 445542 86058 445574 86614
rect 444954 50614 445574 86058
rect 448674 90334 449294 125778
rect 448674 89778 448706 90334
rect 449262 89778 449294 90334
rect 446288 75454 446608 75486
rect 446288 75218 446330 75454
rect 446566 75218 446608 75454
rect 446288 75134 446608 75218
rect 446288 74898 446330 75134
rect 446566 74898 446608 75134
rect 446288 74866 446608 74898
rect 444954 50058 444986 50614
rect 445542 50058 445574 50614
rect 444954 14614 445574 50058
rect 448674 54334 449294 89778
rect 448674 53778 448706 54334
rect 449262 53778 449294 54334
rect 446288 39454 446608 39486
rect 446288 39218 446330 39454
rect 446566 39218 446608 39454
rect 446288 39134 446608 39218
rect 446288 38898 446330 39134
rect 446566 38898 446608 39134
rect 446288 38866 446608 38898
rect 444954 14058 444986 14614
rect 445542 14058 445574 14614
rect 444954 -3226 445574 14058
rect 444954 -3782 444986 -3226
rect 445542 -3782 445574 -3226
rect 444954 -7654 445574 -3782
rect 448674 18334 449294 53778
rect 448674 17778 448706 18334
rect 449262 17778 449294 18334
rect 448674 -4186 449294 17778
rect 448674 -4742 448706 -4186
rect 449262 -4742 449294 -4186
rect 448674 -7654 449294 -4742
rect 452394 709638 453014 711590
rect 452394 709082 452426 709638
rect 452982 709082 453014 709638
rect 452394 670054 453014 709082
rect 452394 669498 452426 670054
rect 452982 669498 453014 670054
rect 452394 634054 453014 669498
rect 452394 633498 452426 634054
rect 452982 633498 453014 634054
rect 452394 598054 453014 633498
rect 452394 597498 452426 598054
rect 452982 597498 453014 598054
rect 452394 562054 453014 597498
rect 452394 561498 452426 562054
rect 452982 561498 453014 562054
rect 452394 526054 453014 561498
rect 452394 525498 452426 526054
rect 452982 525498 453014 526054
rect 452394 490054 453014 525498
rect 452394 489498 452426 490054
rect 452982 489498 453014 490054
rect 452394 454054 453014 489498
rect 452394 453498 452426 454054
rect 452982 453498 453014 454054
rect 452394 418054 453014 453498
rect 452394 417498 452426 418054
rect 452982 417498 453014 418054
rect 452394 382054 453014 417498
rect 452394 381498 452426 382054
rect 452982 381498 453014 382054
rect 452394 346054 453014 381498
rect 452394 345498 452426 346054
rect 452982 345498 453014 346054
rect 452394 310054 453014 345498
rect 452394 309498 452426 310054
rect 452982 309498 453014 310054
rect 452394 274054 453014 309498
rect 452394 273498 452426 274054
rect 452982 273498 453014 274054
rect 452394 238054 453014 273498
rect 452394 237498 452426 238054
rect 452982 237498 453014 238054
rect 452394 202054 453014 237498
rect 452394 201498 452426 202054
rect 452982 201498 453014 202054
rect 452394 166054 453014 201498
rect 452394 165498 452426 166054
rect 452982 165498 453014 166054
rect 452394 130054 453014 165498
rect 452394 129498 452426 130054
rect 452982 129498 453014 130054
rect 452394 94054 453014 129498
rect 452394 93498 452426 94054
rect 452982 93498 453014 94054
rect 452394 58054 453014 93498
rect 452394 57498 452426 58054
rect 452982 57498 453014 58054
rect 452394 22054 453014 57498
rect 452394 21498 452426 22054
rect 452982 21498 453014 22054
rect 452394 -5146 453014 21498
rect 452394 -5702 452426 -5146
rect 452982 -5702 453014 -5146
rect 452394 -7654 453014 -5702
rect 456114 710598 456734 711590
rect 456114 710042 456146 710598
rect 456702 710042 456734 710598
rect 456114 673774 456734 710042
rect 456114 673218 456146 673774
rect 456702 673218 456734 673774
rect 456114 637774 456734 673218
rect 456114 637218 456146 637774
rect 456702 637218 456734 637774
rect 456114 601774 456734 637218
rect 456114 601218 456146 601774
rect 456702 601218 456734 601774
rect 456114 565774 456734 601218
rect 456114 565218 456146 565774
rect 456702 565218 456734 565774
rect 456114 529774 456734 565218
rect 456114 529218 456146 529774
rect 456702 529218 456734 529774
rect 456114 493774 456734 529218
rect 456114 493218 456146 493774
rect 456702 493218 456734 493774
rect 456114 457774 456734 493218
rect 456114 457218 456146 457774
rect 456702 457218 456734 457774
rect 456114 421774 456734 457218
rect 456114 421218 456146 421774
rect 456702 421218 456734 421774
rect 456114 385774 456734 421218
rect 456114 385218 456146 385774
rect 456702 385218 456734 385774
rect 456114 349774 456734 385218
rect 456114 349218 456146 349774
rect 456702 349218 456734 349774
rect 456114 313774 456734 349218
rect 456114 313218 456146 313774
rect 456702 313218 456734 313774
rect 456114 277774 456734 313218
rect 456114 277218 456146 277774
rect 456702 277218 456734 277774
rect 456114 241774 456734 277218
rect 456114 241218 456146 241774
rect 456702 241218 456734 241774
rect 456114 205774 456734 241218
rect 456114 205218 456146 205774
rect 456702 205218 456734 205774
rect 456114 169774 456734 205218
rect 456114 169218 456146 169774
rect 456702 169218 456734 169774
rect 456114 133774 456734 169218
rect 456114 133218 456146 133774
rect 456702 133218 456734 133774
rect 456114 97774 456734 133218
rect 456114 97218 456146 97774
rect 456702 97218 456734 97774
rect 456114 61774 456734 97218
rect 456114 61218 456146 61774
rect 456702 61218 456734 61774
rect 456114 25774 456734 61218
rect 456114 25218 456146 25774
rect 456702 25218 456734 25774
rect 456114 -6106 456734 25218
rect 459834 711558 460454 711590
rect 459834 711002 459866 711558
rect 460422 711002 460454 711558
rect 459834 677494 460454 711002
rect 459834 676938 459866 677494
rect 460422 676938 460454 677494
rect 459834 641494 460454 676938
rect 459834 640938 459866 641494
rect 460422 640938 460454 641494
rect 459834 605494 460454 640938
rect 459834 604938 459866 605494
rect 460422 604938 460454 605494
rect 459834 569494 460454 604938
rect 459834 568938 459866 569494
rect 460422 568938 460454 569494
rect 459834 533494 460454 568938
rect 459834 532938 459866 533494
rect 460422 532938 460454 533494
rect 459834 497494 460454 532938
rect 459834 496938 459866 497494
rect 460422 496938 460454 497494
rect 459834 461494 460454 496938
rect 459834 460938 459866 461494
rect 460422 460938 460454 461494
rect 459834 425494 460454 460938
rect 459834 424938 459866 425494
rect 460422 424938 460454 425494
rect 459834 389494 460454 424938
rect 459834 388938 459866 389494
rect 460422 388938 460454 389494
rect 459834 353494 460454 388938
rect 459834 352938 459866 353494
rect 460422 352938 460454 353494
rect 459834 317494 460454 352938
rect 469794 704838 470414 711590
rect 469794 704282 469826 704838
rect 470382 704282 470414 704838
rect 469794 687454 470414 704282
rect 469794 686898 469826 687454
rect 470382 686898 470414 687454
rect 469794 651454 470414 686898
rect 469794 650898 469826 651454
rect 470382 650898 470414 651454
rect 469794 615454 470414 650898
rect 469794 614898 469826 615454
rect 470382 614898 470414 615454
rect 469794 579454 470414 614898
rect 469794 578898 469826 579454
rect 470382 578898 470414 579454
rect 469794 543454 470414 578898
rect 469794 542898 469826 543454
rect 470382 542898 470414 543454
rect 469794 507454 470414 542898
rect 469794 506898 469826 507454
rect 470382 506898 470414 507454
rect 469794 471454 470414 506898
rect 469794 470898 469826 471454
rect 470382 470898 470414 471454
rect 469794 435454 470414 470898
rect 469794 434898 469826 435454
rect 470382 434898 470414 435454
rect 469794 399454 470414 434898
rect 469794 398898 469826 399454
rect 470382 398898 470414 399454
rect 469794 363454 470414 398898
rect 469794 362898 469826 363454
rect 470382 362898 470414 363454
rect 461648 331174 461968 331206
rect 461648 330938 461690 331174
rect 461926 330938 461968 331174
rect 461648 330854 461968 330938
rect 461648 330618 461690 330854
rect 461926 330618 461968 330854
rect 461648 330586 461968 330618
rect 459834 316938 459866 317494
rect 460422 316938 460454 317494
rect 459834 281494 460454 316938
rect 469794 327454 470414 362898
rect 469794 326898 469826 327454
rect 470382 326898 470414 327454
rect 461648 295174 461968 295206
rect 461648 294938 461690 295174
rect 461926 294938 461968 295174
rect 461648 294854 461968 294938
rect 461648 294618 461690 294854
rect 461926 294618 461968 294854
rect 461648 294586 461968 294618
rect 459834 280938 459866 281494
rect 460422 280938 460454 281494
rect 459834 245494 460454 280938
rect 469794 291454 470414 326898
rect 469794 290898 469826 291454
rect 470382 290898 470414 291454
rect 461648 259174 461968 259206
rect 461648 258938 461690 259174
rect 461926 258938 461968 259174
rect 461648 258854 461968 258938
rect 461648 258618 461690 258854
rect 461926 258618 461968 258854
rect 461648 258586 461968 258618
rect 459834 244938 459866 245494
rect 460422 244938 460454 245494
rect 459834 209494 460454 244938
rect 469794 255454 470414 290898
rect 469794 254898 469826 255454
rect 470382 254898 470414 255454
rect 461648 223174 461968 223206
rect 461648 222938 461690 223174
rect 461926 222938 461968 223174
rect 461648 222854 461968 222938
rect 461648 222618 461690 222854
rect 461926 222618 461968 222854
rect 461648 222586 461968 222618
rect 459834 208938 459866 209494
rect 460422 208938 460454 209494
rect 459834 173494 460454 208938
rect 469794 219454 470414 254898
rect 469794 218898 469826 219454
rect 470382 218898 470414 219454
rect 461648 187174 461968 187206
rect 461648 186938 461690 187174
rect 461926 186938 461968 187174
rect 461648 186854 461968 186938
rect 461648 186618 461690 186854
rect 461926 186618 461968 186854
rect 461648 186586 461968 186618
rect 459834 172938 459866 173494
rect 460422 172938 460454 173494
rect 459834 137494 460454 172938
rect 469794 183454 470414 218898
rect 469794 182898 469826 183454
rect 470382 182898 470414 183454
rect 461648 151174 461968 151206
rect 461648 150938 461690 151174
rect 461926 150938 461968 151174
rect 461648 150854 461968 150938
rect 461648 150618 461690 150854
rect 461926 150618 461968 150854
rect 461648 150586 461968 150618
rect 459834 136938 459866 137494
rect 460422 136938 460454 137494
rect 459834 101494 460454 136938
rect 469794 147454 470414 182898
rect 469794 146898 469826 147454
rect 470382 146898 470414 147454
rect 461648 115174 461968 115206
rect 461648 114938 461690 115174
rect 461926 114938 461968 115174
rect 461648 114854 461968 114938
rect 461648 114618 461690 114854
rect 461926 114618 461968 114854
rect 461648 114586 461968 114618
rect 459834 100938 459866 101494
rect 460422 100938 460454 101494
rect 459834 65494 460454 100938
rect 469794 111454 470414 146898
rect 469794 110898 469826 111454
rect 470382 110898 470414 111454
rect 461648 79174 461968 79206
rect 461648 78938 461690 79174
rect 461926 78938 461968 79174
rect 461648 78854 461968 78938
rect 461648 78618 461690 78854
rect 461926 78618 461968 78854
rect 461648 78586 461968 78618
rect 459834 64938 459866 65494
rect 460422 64938 460454 65494
rect 459834 29494 460454 64938
rect 469794 75454 470414 110898
rect 469794 74898 469826 75454
rect 470382 74898 470414 75454
rect 461648 43174 461968 43206
rect 461648 42938 461690 43174
rect 461926 42938 461968 43174
rect 461648 42854 461968 42938
rect 461648 42618 461690 42854
rect 461926 42618 461968 42854
rect 461648 42586 461968 42618
rect 459834 28938 459866 29494
rect 460422 28938 460454 29494
rect 458403 3364 458469 3365
rect 458403 3300 458404 3364
rect 458468 3300 458469 3364
rect 458403 3299 458469 3300
rect 458406 2957 458466 3299
rect 458403 2956 458469 2957
rect 458403 2892 458404 2956
rect 458468 2892 458469 2956
rect 458403 2891 458469 2892
rect 456114 -6662 456146 -6106
rect 456702 -6662 456734 -6106
rect 456114 -7654 456734 -6662
rect 459834 -7066 460454 28938
rect 469794 39454 470414 74898
rect 469794 38898 469826 39454
rect 470382 38898 470414 39454
rect 461648 7174 461968 7206
rect 461648 6938 461690 7174
rect 461926 6938 461968 7174
rect 461648 6854 461968 6938
rect 461648 6618 461690 6854
rect 461926 6618 461968 6854
rect 461648 6586 461968 6618
rect 462635 3636 462701 3637
rect 462635 3572 462636 3636
rect 462700 3572 462701 3636
rect 462635 3571 462701 3572
rect 462638 2685 462698 3571
rect 463739 3500 463805 3501
rect 463739 3436 463740 3500
rect 463804 3436 463805 3500
rect 463739 3435 463805 3436
rect 469794 3454 470414 38898
rect 463742 2821 463802 3435
rect 467235 3364 467301 3365
rect 467235 3300 467236 3364
rect 467300 3300 467301 3364
rect 467235 3299 467301 3300
rect 466315 3228 466381 3229
rect 466315 3164 466316 3228
rect 466380 3164 466381 3228
rect 466315 3163 466381 3164
rect 463739 2820 463805 2821
rect 463739 2756 463740 2820
rect 463804 2756 463805 2820
rect 463739 2755 463805 2756
rect 462635 2684 462701 2685
rect 462635 2620 462636 2684
rect 462700 2620 462701 2684
rect 462635 2619 462701 2620
rect 466318 2549 466378 3163
rect 467238 2549 467298 3299
rect 469794 2898 469826 3454
rect 470382 2898 470414 3454
rect 466315 2548 466381 2549
rect 466315 2484 466316 2548
rect 466380 2484 466381 2548
rect 466315 2483 466381 2484
rect 467235 2548 467301 2549
rect 467235 2484 467236 2548
rect 467300 2484 467301 2548
rect 467235 2483 467301 2484
rect 459834 -7622 459866 -7066
rect 460422 -7622 460454 -7066
rect 459834 -7654 460454 -7622
rect 469794 -346 470414 2898
rect 469794 -902 469826 -346
rect 470382 -902 470414 -346
rect 469794 -7654 470414 -902
rect 473514 705798 474134 711590
rect 473514 705242 473546 705798
rect 474102 705242 474134 705798
rect 473514 691174 474134 705242
rect 473514 690618 473546 691174
rect 474102 690618 474134 691174
rect 473514 655174 474134 690618
rect 473514 654618 473546 655174
rect 474102 654618 474134 655174
rect 473514 619174 474134 654618
rect 473514 618618 473546 619174
rect 474102 618618 474134 619174
rect 473514 583174 474134 618618
rect 473514 582618 473546 583174
rect 474102 582618 474134 583174
rect 473514 547174 474134 582618
rect 473514 546618 473546 547174
rect 474102 546618 474134 547174
rect 473514 511174 474134 546618
rect 473514 510618 473546 511174
rect 474102 510618 474134 511174
rect 473514 475174 474134 510618
rect 473514 474618 473546 475174
rect 474102 474618 474134 475174
rect 473514 439174 474134 474618
rect 473514 438618 473546 439174
rect 474102 438618 474134 439174
rect 473514 403174 474134 438618
rect 473514 402618 473546 403174
rect 474102 402618 474134 403174
rect 473514 367174 474134 402618
rect 473514 366618 473546 367174
rect 474102 366618 474134 367174
rect 473514 331174 474134 366618
rect 477234 706758 477854 711590
rect 477234 706202 477266 706758
rect 477822 706202 477854 706758
rect 477234 694894 477854 706202
rect 477234 694338 477266 694894
rect 477822 694338 477854 694894
rect 477234 658894 477854 694338
rect 477234 658338 477266 658894
rect 477822 658338 477854 658894
rect 477234 622894 477854 658338
rect 477234 622338 477266 622894
rect 477822 622338 477854 622894
rect 477234 586894 477854 622338
rect 477234 586338 477266 586894
rect 477822 586338 477854 586894
rect 477234 550894 477854 586338
rect 477234 550338 477266 550894
rect 477822 550338 477854 550894
rect 477234 514894 477854 550338
rect 477234 514338 477266 514894
rect 477822 514338 477854 514894
rect 477234 478894 477854 514338
rect 477234 478338 477266 478894
rect 477822 478338 477854 478894
rect 477234 442894 477854 478338
rect 477234 442338 477266 442894
rect 477822 442338 477854 442894
rect 477234 406894 477854 442338
rect 477234 406338 477266 406894
rect 477822 406338 477854 406894
rect 477234 370894 477854 406338
rect 477234 370338 477266 370894
rect 477822 370338 477854 370894
rect 477234 354980 477854 370338
rect 480954 707718 481574 711590
rect 480954 707162 480986 707718
rect 481542 707162 481574 707718
rect 480954 698614 481574 707162
rect 480954 698058 480986 698614
rect 481542 698058 481574 698614
rect 480954 662614 481574 698058
rect 480954 662058 480986 662614
rect 481542 662058 481574 662614
rect 480954 626614 481574 662058
rect 480954 626058 480986 626614
rect 481542 626058 481574 626614
rect 480954 590614 481574 626058
rect 480954 590058 480986 590614
rect 481542 590058 481574 590614
rect 480954 554614 481574 590058
rect 480954 554058 480986 554614
rect 481542 554058 481574 554614
rect 480954 518614 481574 554058
rect 480954 518058 480986 518614
rect 481542 518058 481574 518614
rect 480954 482614 481574 518058
rect 480954 482058 480986 482614
rect 481542 482058 481574 482614
rect 480954 446614 481574 482058
rect 480954 446058 480986 446614
rect 481542 446058 481574 446614
rect 480954 410614 481574 446058
rect 480954 410058 480986 410614
rect 481542 410058 481574 410614
rect 480954 374614 481574 410058
rect 480954 374058 480986 374614
rect 481542 374058 481574 374614
rect 473514 330618 473546 331174
rect 474102 330618 474134 331174
rect 473514 295174 474134 330618
rect 480954 338614 481574 374058
rect 480954 338058 480986 338614
rect 481542 338058 481574 338614
rect 477008 327454 477328 327486
rect 477008 327218 477050 327454
rect 477286 327218 477328 327454
rect 477008 327134 477328 327218
rect 477008 326898 477050 327134
rect 477286 326898 477328 327134
rect 477008 326866 477328 326898
rect 473514 294618 473546 295174
rect 474102 294618 474134 295174
rect 473514 259174 474134 294618
rect 480954 302614 481574 338058
rect 480954 302058 480986 302614
rect 481542 302058 481574 302614
rect 477008 291454 477328 291486
rect 477008 291218 477050 291454
rect 477286 291218 477328 291454
rect 477008 291134 477328 291218
rect 477008 290898 477050 291134
rect 477286 290898 477328 291134
rect 477008 290866 477328 290898
rect 473514 258618 473546 259174
rect 474102 258618 474134 259174
rect 473514 223174 474134 258618
rect 480954 266614 481574 302058
rect 480954 266058 480986 266614
rect 481542 266058 481574 266614
rect 477008 255454 477328 255486
rect 477008 255218 477050 255454
rect 477286 255218 477328 255454
rect 477008 255134 477328 255218
rect 477008 254898 477050 255134
rect 477286 254898 477328 255134
rect 477008 254866 477328 254898
rect 473514 222618 473546 223174
rect 474102 222618 474134 223174
rect 473514 187174 474134 222618
rect 480954 230614 481574 266058
rect 480954 230058 480986 230614
rect 481542 230058 481574 230614
rect 477008 219454 477328 219486
rect 477008 219218 477050 219454
rect 477286 219218 477328 219454
rect 477008 219134 477328 219218
rect 477008 218898 477050 219134
rect 477286 218898 477328 219134
rect 477008 218866 477328 218898
rect 473514 186618 473546 187174
rect 474102 186618 474134 187174
rect 473514 151174 474134 186618
rect 480954 194614 481574 230058
rect 480954 194058 480986 194614
rect 481542 194058 481574 194614
rect 477008 183454 477328 183486
rect 477008 183218 477050 183454
rect 477286 183218 477328 183454
rect 477008 183134 477328 183218
rect 477008 182898 477050 183134
rect 477286 182898 477328 183134
rect 477008 182866 477328 182898
rect 473514 150618 473546 151174
rect 474102 150618 474134 151174
rect 473514 115174 474134 150618
rect 480954 158614 481574 194058
rect 480954 158058 480986 158614
rect 481542 158058 481574 158614
rect 477008 147454 477328 147486
rect 477008 147218 477050 147454
rect 477286 147218 477328 147454
rect 477008 147134 477328 147218
rect 477008 146898 477050 147134
rect 477286 146898 477328 147134
rect 477008 146866 477328 146898
rect 473514 114618 473546 115174
rect 474102 114618 474134 115174
rect 473514 79174 474134 114618
rect 480954 122614 481574 158058
rect 480954 122058 480986 122614
rect 481542 122058 481574 122614
rect 477008 111454 477328 111486
rect 477008 111218 477050 111454
rect 477286 111218 477328 111454
rect 477008 111134 477328 111218
rect 477008 110898 477050 111134
rect 477286 110898 477328 111134
rect 477008 110866 477328 110898
rect 473514 78618 473546 79174
rect 474102 78618 474134 79174
rect 473514 43174 474134 78618
rect 480954 86614 481574 122058
rect 480954 86058 480986 86614
rect 481542 86058 481574 86614
rect 477008 75454 477328 75486
rect 477008 75218 477050 75454
rect 477286 75218 477328 75454
rect 477008 75134 477328 75218
rect 477008 74898 477050 75134
rect 477286 74898 477328 75134
rect 477008 74866 477328 74898
rect 473514 42618 473546 43174
rect 474102 42618 474134 43174
rect 473514 7174 474134 42618
rect 480954 50614 481574 86058
rect 480954 50058 480986 50614
rect 481542 50058 481574 50614
rect 477008 39454 477328 39486
rect 477008 39218 477050 39454
rect 477286 39218 477328 39454
rect 477008 39134 477328 39218
rect 477008 38898 477050 39134
rect 477286 38898 477328 39134
rect 477008 38866 477328 38898
rect 473514 6618 473546 7174
rect 474102 6618 474134 7174
rect 473514 -1306 474134 6618
rect 473514 -1862 473546 -1306
rect 474102 -1862 474134 -1306
rect 473514 -7654 474134 -1862
rect 480954 14614 481574 50058
rect 480954 14058 480986 14614
rect 481542 14058 481574 14614
rect 480954 -3226 481574 14058
rect 480954 -3782 480986 -3226
rect 481542 -3782 481574 -3226
rect 480954 -7654 481574 -3782
rect 484674 708678 485294 711590
rect 484674 708122 484706 708678
rect 485262 708122 485294 708678
rect 484674 666334 485294 708122
rect 484674 665778 484706 666334
rect 485262 665778 485294 666334
rect 484674 630334 485294 665778
rect 484674 629778 484706 630334
rect 485262 629778 485294 630334
rect 484674 594334 485294 629778
rect 484674 593778 484706 594334
rect 485262 593778 485294 594334
rect 484674 558334 485294 593778
rect 484674 557778 484706 558334
rect 485262 557778 485294 558334
rect 484674 522334 485294 557778
rect 484674 521778 484706 522334
rect 485262 521778 485294 522334
rect 484674 486334 485294 521778
rect 484674 485778 484706 486334
rect 485262 485778 485294 486334
rect 484674 450334 485294 485778
rect 484674 449778 484706 450334
rect 485262 449778 485294 450334
rect 484674 414334 485294 449778
rect 484674 413778 484706 414334
rect 485262 413778 485294 414334
rect 484674 378334 485294 413778
rect 484674 377778 484706 378334
rect 485262 377778 485294 378334
rect 484674 342334 485294 377778
rect 484674 341778 484706 342334
rect 485262 341778 485294 342334
rect 484674 306334 485294 341778
rect 484674 305778 484706 306334
rect 485262 305778 485294 306334
rect 484674 270334 485294 305778
rect 484674 269778 484706 270334
rect 485262 269778 485294 270334
rect 484674 234334 485294 269778
rect 484674 233778 484706 234334
rect 485262 233778 485294 234334
rect 484674 198334 485294 233778
rect 484674 197778 484706 198334
rect 485262 197778 485294 198334
rect 484674 162334 485294 197778
rect 484674 161778 484706 162334
rect 485262 161778 485294 162334
rect 484674 126334 485294 161778
rect 484674 125778 484706 126334
rect 485262 125778 485294 126334
rect 484674 90334 485294 125778
rect 484674 89778 484706 90334
rect 485262 89778 485294 90334
rect 484674 54334 485294 89778
rect 484674 53778 484706 54334
rect 485262 53778 485294 54334
rect 484674 18334 485294 53778
rect 484674 17778 484706 18334
rect 485262 17778 485294 18334
rect 484674 -4186 485294 17778
rect 484674 -4742 484706 -4186
rect 485262 -4742 485294 -4186
rect 484674 -7654 485294 -4742
rect 488394 709638 489014 711590
rect 488394 709082 488426 709638
rect 488982 709082 489014 709638
rect 488394 670054 489014 709082
rect 488394 669498 488426 670054
rect 488982 669498 489014 670054
rect 488394 634054 489014 669498
rect 488394 633498 488426 634054
rect 488982 633498 489014 634054
rect 488394 598054 489014 633498
rect 488394 597498 488426 598054
rect 488982 597498 489014 598054
rect 488394 562054 489014 597498
rect 488394 561498 488426 562054
rect 488982 561498 489014 562054
rect 488394 526054 489014 561498
rect 488394 525498 488426 526054
rect 488982 525498 489014 526054
rect 488394 490054 489014 525498
rect 488394 489498 488426 490054
rect 488982 489498 489014 490054
rect 488394 454054 489014 489498
rect 488394 453498 488426 454054
rect 488982 453498 489014 454054
rect 488394 418054 489014 453498
rect 488394 417498 488426 418054
rect 488982 417498 489014 418054
rect 488394 382054 489014 417498
rect 488394 381498 488426 382054
rect 488982 381498 489014 382054
rect 488394 346054 489014 381498
rect 492114 710598 492734 711590
rect 492114 710042 492146 710598
rect 492702 710042 492734 710598
rect 492114 673774 492734 710042
rect 492114 673218 492146 673774
rect 492702 673218 492734 673774
rect 492114 637774 492734 673218
rect 492114 637218 492146 637774
rect 492702 637218 492734 637774
rect 492114 601774 492734 637218
rect 492114 601218 492146 601774
rect 492702 601218 492734 601774
rect 492114 565774 492734 601218
rect 492114 565218 492146 565774
rect 492702 565218 492734 565774
rect 492114 529774 492734 565218
rect 492114 529218 492146 529774
rect 492702 529218 492734 529774
rect 492114 493774 492734 529218
rect 492114 493218 492146 493774
rect 492702 493218 492734 493774
rect 492114 457774 492734 493218
rect 492114 457218 492146 457774
rect 492702 457218 492734 457774
rect 492114 421774 492734 457218
rect 492114 421218 492146 421774
rect 492702 421218 492734 421774
rect 492114 385774 492734 421218
rect 492114 385218 492146 385774
rect 492702 385218 492734 385774
rect 492114 354980 492734 385218
rect 495834 711558 496454 711590
rect 495834 711002 495866 711558
rect 496422 711002 496454 711558
rect 495834 677494 496454 711002
rect 495834 676938 495866 677494
rect 496422 676938 496454 677494
rect 495834 641494 496454 676938
rect 495834 640938 495866 641494
rect 496422 640938 496454 641494
rect 495834 605494 496454 640938
rect 495834 604938 495866 605494
rect 496422 604938 496454 605494
rect 495834 569494 496454 604938
rect 495834 568938 495866 569494
rect 496422 568938 496454 569494
rect 495834 533494 496454 568938
rect 495834 532938 495866 533494
rect 496422 532938 496454 533494
rect 495834 497494 496454 532938
rect 495834 496938 495866 497494
rect 496422 496938 496454 497494
rect 495834 461494 496454 496938
rect 495834 460938 495866 461494
rect 496422 460938 496454 461494
rect 495834 425494 496454 460938
rect 495834 424938 495866 425494
rect 496422 424938 496454 425494
rect 495834 389494 496454 424938
rect 495834 388938 495866 389494
rect 496422 388938 496454 389494
rect 488394 345498 488426 346054
rect 488982 345498 489014 346054
rect 488394 310054 489014 345498
rect 495834 353494 496454 388938
rect 495834 352938 495866 353494
rect 496422 352938 496454 353494
rect 492368 331174 492688 331206
rect 492368 330938 492410 331174
rect 492646 330938 492688 331174
rect 492368 330854 492688 330938
rect 492368 330618 492410 330854
rect 492646 330618 492688 330854
rect 492368 330586 492688 330618
rect 488394 309498 488426 310054
rect 488982 309498 489014 310054
rect 488394 274054 489014 309498
rect 495834 317494 496454 352938
rect 495834 316938 495866 317494
rect 496422 316938 496454 317494
rect 492368 295174 492688 295206
rect 492368 294938 492410 295174
rect 492646 294938 492688 295174
rect 492368 294854 492688 294938
rect 492368 294618 492410 294854
rect 492646 294618 492688 294854
rect 492368 294586 492688 294618
rect 488394 273498 488426 274054
rect 488982 273498 489014 274054
rect 488394 238054 489014 273498
rect 495834 281494 496454 316938
rect 495834 280938 495866 281494
rect 496422 280938 496454 281494
rect 492368 259174 492688 259206
rect 492368 258938 492410 259174
rect 492646 258938 492688 259174
rect 492368 258854 492688 258938
rect 492368 258618 492410 258854
rect 492646 258618 492688 258854
rect 492368 258586 492688 258618
rect 488394 237498 488426 238054
rect 488982 237498 489014 238054
rect 488394 202054 489014 237498
rect 495834 245494 496454 280938
rect 495834 244938 495866 245494
rect 496422 244938 496454 245494
rect 492368 223174 492688 223206
rect 492368 222938 492410 223174
rect 492646 222938 492688 223174
rect 492368 222854 492688 222938
rect 492368 222618 492410 222854
rect 492646 222618 492688 222854
rect 492368 222586 492688 222618
rect 488394 201498 488426 202054
rect 488982 201498 489014 202054
rect 488394 166054 489014 201498
rect 495834 209494 496454 244938
rect 495834 208938 495866 209494
rect 496422 208938 496454 209494
rect 492368 187174 492688 187206
rect 492368 186938 492410 187174
rect 492646 186938 492688 187174
rect 492368 186854 492688 186938
rect 492368 186618 492410 186854
rect 492646 186618 492688 186854
rect 492368 186586 492688 186618
rect 488394 165498 488426 166054
rect 488982 165498 489014 166054
rect 488394 130054 489014 165498
rect 495834 173494 496454 208938
rect 495834 172938 495866 173494
rect 496422 172938 496454 173494
rect 492368 151174 492688 151206
rect 492368 150938 492410 151174
rect 492646 150938 492688 151174
rect 492368 150854 492688 150938
rect 492368 150618 492410 150854
rect 492646 150618 492688 150854
rect 492368 150586 492688 150618
rect 488394 129498 488426 130054
rect 488982 129498 489014 130054
rect 488394 94054 489014 129498
rect 495834 137494 496454 172938
rect 495834 136938 495866 137494
rect 496422 136938 496454 137494
rect 492368 115174 492688 115206
rect 492368 114938 492410 115174
rect 492646 114938 492688 115174
rect 492368 114854 492688 114938
rect 492368 114618 492410 114854
rect 492646 114618 492688 114854
rect 492368 114586 492688 114618
rect 488394 93498 488426 94054
rect 488982 93498 489014 94054
rect 488394 58054 489014 93498
rect 495834 101494 496454 136938
rect 495834 100938 495866 101494
rect 496422 100938 496454 101494
rect 492368 79174 492688 79206
rect 492368 78938 492410 79174
rect 492646 78938 492688 79174
rect 492368 78854 492688 78938
rect 492368 78618 492410 78854
rect 492646 78618 492688 78854
rect 492368 78586 492688 78618
rect 488394 57498 488426 58054
rect 488982 57498 489014 58054
rect 488394 22054 489014 57498
rect 495834 65494 496454 100938
rect 495834 64938 495866 65494
rect 496422 64938 496454 65494
rect 492368 43174 492688 43206
rect 492368 42938 492410 43174
rect 492646 42938 492688 43174
rect 492368 42854 492688 42938
rect 492368 42618 492410 42854
rect 492646 42618 492688 42854
rect 492368 42586 492688 42618
rect 488394 21498 488426 22054
rect 488982 21498 489014 22054
rect 488394 -5146 489014 21498
rect 495834 29494 496454 64938
rect 495834 28938 495866 29494
rect 496422 28938 496454 29494
rect 492368 7174 492688 7206
rect 492368 6938 492410 7174
rect 492646 6938 492688 7174
rect 492368 6854 492688 6938
rect 492368 6618 492410 6854
rect 492646 6618 492688 6854
rect 492368 6586 492688 6618
rect 488394 -5702 488426 -5146
rect 488982 -5702 489014 -5146
rect 488394 -7654 489014 -5702
rect 495834 -7066 496454 28938
rect 505794 704838 506414 711590
rect 505794 704282 505826 704838
rect 506382 704282 506414 704838
rect 505794 687454 506414 704282
rect 505794 686898 505826 687454
rect 506382 686898 506414 687454
rect 505794 651454 506414 686898
rect 505794 650898 505826 651454
rect 506382 650898 506414 651454
rect 505794 615454 506414 650898
rect 505794 614898 505826 615454
rect 506382 614898 506414 615454
rect 505794 579454 506414 614898
rect 505794 578898 505826 579454
rect 506382 578898 506414 579454
rect 505794 543454 506414 578898
rect 505794 542898 505826 543454
rect 506382 542898 506414 543454
rect 505794 507454 506414 542898
rect 505794 506898 505826 507454
rect 506382 506898 506414 507454
rect 505794 471454 506414 506898
rect 505794 470898 505826 471454
rect 506382 470898 506414 471454
rect 505794 435454 506414 470898
rect 505794 434898 505826 435454
rect 506382 434898 506414 435454
rect 505794 399454 506414 434898
rect 505794 398898 505826 399454
rect 506382 398898 506414 399454
rect 505794 363454 506414 398898
rect 505794 362898 505826 363454
rect 506382 362898 506414 363454
rect 505794 327454 506414 362898
rect 509514 705798 510134 711590
rect 509514 705242 509546 705798
rect 510102 705242 510134 705798
rect 509514 691174 510134 705242
rect 509514 690618 509546 691174
rect 510102 690618 510134 691174
rect 509514 655174 510134 690618
rect 509514 654618 509546 655174
rect 510102 654618 510134 655174
rect 509514 619174 510134 654618
rect 509514 618618 509546 619174
rect 510102 618618 510134 619174
rect 509514 583174 510134 618618
rect 509514 582618 509546 583174
rect 510102 582618 510134 583174
rect 509514 547174 510134 582618
rect 509514 546618 509546 547174
rect 510102 546618 510134 547174
rect 509514 511174 510134 546618
rect 509514 510618 509546 511174
rect 510102 510618 510134 511174
rect 509514 475174 510134 510618
rect 509514 474618 509546 475174
rect 510102 474618 510134 475174
rect 509514 439174 510134 474618
rect 509514 438618 509546 439174
rect 510102 438618 510134 439174
rect 509514 403174 510134 438618
rect 509514 402618 509546 403174
rect 510102 402618 510134 403174
rect 509514 367174 510134 402618
rect 509514 366618 509546 367174
rect 510102 366618 510134 367174
rect 509514 331174 510134 366618
rect 509514 330618 509546 331174
rect 510102 330618 510134 331174
rect 505794 326898 505826 327454
rect 506382 326898 506414 327454
rect 505794 291454 506414 326898
rect 507728 327454 508048 327486
rect 507728 327218 507770 327454
rect 508006 327218 508048 327454
rect 507728 327134 508048 327218
rect 507728 326898 507770 327134
rect 508006 326898 508048 327134
rect 507728 326866 508048 326898
rect 509514 295174 510134 330618
rect 509514 294618 509546 295174
rect 510102 294618 510134 295174
rect 505794 290898 505826 291454
rect 506382 290898 506414 291454
rect 505794 255454 506414 290898
rect 507728 291454 508048 291486
rect 507728 291218 507770 291454
rect 508006 291218 508048 291454
rect 507728 291134 508048 291218
rect 507728 290898 507770 291134
rect 508006 290898 508048 291134
rect 507728 290866 508048 290898
rect 509514 259174 510134 294618
rect 509514 258618 509546 259174
rect 510102 258618 510134 259174
rect 505794 254898 505826 255454
rect 506382 254898 506414 255454
rect 505794 219454 506414 254898
rect 507728 255454 508048 255486
rect 507728 255218 507770 255454
rect 508006 255218 508048 255454
rect 507728 255134 508048 255218
rect 507728 254898 507770 255134
rect 508006 254898 508048 255134
rect 507728 254866 508048 254898
rect 509514 223174 510134 258618
rect 509514 222618 509546 223174
rect 510102 222618 510134 223174
rect 505794 218898 505826 219454
rect 506382 218898 506414 219454
rect 505794 183454 506414 218898
rect 507728 219454 508048 219486
rect 507728 219218 507770 219454
rect 508006 219218 508048 219454
rect 507728 219134 508048 219218
rect 507728 218898 507770 219134
rect 508006 218898 508048 219134
rect 507728 218866 508048 218898
rect 509514 187174 510134 222618
rect 509514 186618 509546 187174
rect 510102 186618 510134 187174
rect 505794 182898 505826 183454
rect 506382 182898 506414 183454
rect 505794 147454 506414 182898
rect 507728 183454 508048 183486
rect 507728 183218 507770 183454
rect 508006 183218 508048 183454
rect 507728 183134 508048 183218
rect 507728 182898 507770 183134
rect 508006 182898 508048 183134
rect 507728 182866 508048 182898
rect 509514 151174 510134 186618
rect 509514 150618 509546 151174
rect 510102 150618 510134 151174
rect 505794 146898 505826 147454
rect 506382 146898 506414 147454
rect 505794 111454 506414 146898
rect 507728 147454 508048 147486
rect 507728 147218 507770 147454
rect 508006 147218 508048 147454
rect 507728 147134 508048 147218
rect 507728 146898 507770 147134
rect 508006 146898 508048 147134
rect 507728 146866 508048 146898
rect 509514 115174 510134 150618
rect 509514 114618 509546 115174
rect 510102 114618 510134 115174
rect 505794 110898 505826 111454
rect 506382 110898 506414 111454
rect 505794 75454 506414 110898
rect 507728 111454 508048 111486
rect 507728 111218 507770 111454
rect 508006 111218 508048 111454
rect 507728 111134 508048 111218
rect 507728 110898 507770 111134
rect 508006 110898 508048 111134
rect 507728 110866 508048 110898
rect 509514 79174 510134 114618
rect 509514 78618 509546 79174
rect 510102 78618 510134 79174
rect 505794 74898 505826 75454
rect 506382 74898 506414 75454
rect 505794 39454 506414 74898
rect 507728 75454 508048 75486
rect 507728 75218 507770 75454
rect 508006 75218 508048 75454
rect 507728 75134 508048 75218
rect 507728 74898 507770 75134
rect 508006 74898 508048 75134
rect 507728 74866 508048 74898
rect 509514 43174 510134 78618
rect 509514 42618 509546 43174
rect 510102 42618 510134 43174
rect 505794 38898 505826 39454
rect 506382 38898 506414 39454
rect 505794 3454 506414 38898
rect 507728 39454 508048 39486
rect 507728 39218 507770 39454
rect 508006 39218 508048 39454
rect 507728 39134 508048 39218
rect 507728 38898 507770 39134
rect 508006 38898 508048 39134
rect 507728 38866 508048 38898
rect 498147 3092 498213 3093
rect 498147 3028 498148 3092
rect 498212 3028 498213 3092
rect 498147 3027 498213 3028
rect 498150 2549 498210 3027
rect 505794 2898 505826 3454
rect 506382 2898 506414 3454
rect 498147 2548 498213 2549
rect 498147 2484 498148 2548
rect 498212 2484 498213 2548
rect 498147 2483 498213 2484
rect 495834 -7622 495866 -7066
rect 496422 -7622 496454 -7066
rect 495834 -7654 496454 -7622
rect 505794 -346 506414 2898
rect 505794 -902 505826 -346
rect 506382 -902 506414 -346
rect 505794 -7654 506414 -902
rect 509514 7174 510134 42618
rect 509514 6618 509546 7174
rect 510102 6618 510134 7174
rect 509514 -1306 510134 6618
rect 509514 -1862 509546 -1306
rect 510102 -1862 510134 -1306
rect 509514 -7654 510134 -1862
rect 513234 706758 513854 711590
rect 513234 706202 513266 706758
rect 513822 706202 513854 706758
rect 513234 694894 513854 706202
rect 513234 694338 513266 694894
rect 513822 694338 513854 694894
rect 513234 658894 513854 694338
rect 513234 658338 513266 658894
rect 513822 658338 513854 658894
rect 513234 622894 513854 658338
rect 513234 622338 513266 622894
rect 513822 622338 513854 622894
rect 513234 586894 513854 622338
rect 513234 586338 513266 586894
rect 513822 586338 513854 586894
rect 513234 550894 513854 586338
rect 513234 550338 513266 550894
rect 513822 550338 513854 550894
rect 513234 514894 513854 550338
rect 513234 514338 513266 514894
rect 513822 514338 513854 514894
rect 513234 478894 513854 514338
rect 513234 478338 513266 478894
rect 513822 478338 513854 478894
rect 513234 442894 513854 478338
rect 513234 442338 513266 442894
rect 513822 442338 513854 442894
rect 513234 406894 513854 442338
rect 513234 406338 513266 406894
rect 513822 406338 513854 406894
rect 513234 370894 513854 406338
rect 513234 370338 513266 370894
rect 513822 370338 513854 370894
rect 513234 334894 513854 370338
rect 513234 334338 513266 334894
rect 513822 334338 513854 334894
rect 513234 298894 513854 334338
rect 513234 298338 513266 298894
rect 513822 298338 513854 298894
rect 513234 262894 513854 298338
rect 513234 262338 513266 262894
rect 513822 262338 513854 262894
rect 513234 226894 513854 262338
rect 513234 226338 513266 226894
rect 513822 226338 513854 226894
rect 513234 190894 513854 226338
rect 513234 190338 513266 190894
rect 513822 190338 513854 190894
rect 513234 154894 513854 190338
rect 513234 154338 513266 154894
rect 513822 154338 513854 154894
rect 513234 118894 513854 154338
rect 513234 118338 513266 118894
rect 513822 118338 513854 118894
rect 513234 82894 513854 118338
rect 513234 82338 513266 82894
rect 513822 82338 513854 82894
rect 513234 46894 513854 82338
rect 513234 46338 513266 46894
rect 513822 46338 513854 46894
rect 513234 10894 513854 46338
rect 513234 10338 513266 10894
rect 513822 10338 513854 10894
rect 513234 -2266 513854 10338
rect 516954 707718 517574 711590
rect 516954 707162 516986 707718
rect 517542 707162 517574 707718
rect 516954 698614 517574 707162
rect 516954 698058 516986 698614
rect 517542 698058 517574 698614
rect 516954 662614 517574 698058
rect 516954 662058 516986 662614
rect 517542 662058 517574 662614
rect 516954 626614 517574 662058
rect 516954 626058 516986 626614
rect 517542 626058 517574 626614
rect 516954 590614 517574 626058
rect 516954 590058 516986 590614
rect 517542 590058 517574 590614
rect 516954 554614 517574 590058
rect 516954 554058 516986 554614
rect 517542 554058 517574 554614
rect 516954 518614 517574 554058
rect 516954 518058 516986 518614
rect 517542 518058 517574 518614
rect 516954 482614 517574 518058
rect 516954 482058 516986 482614
rect 517542 482058 517574 482614
rect 516954 446614 517574 482058
rect 516954 446058 516986 446614
rect 517542 446058 517574 446614
rect 516954 410614 517574 446058
rect 516954 410058 516986 410614
rect 517542 410058 517574 410614
rect 516954 374614 517574 410058
rect 516954 374058 516986 374614
rect 517542 374058 517574 374614
rect 516954 338614 517574 374058
rect 516954 338058 516986 338614
rect 517542 338058 517574 338614
rect 516954 302614 517574 338058
rect 516954 302058 516986 302614
rect 517542 302058 517574 302614
rect 516954 266614 517574 302058
rect 516954 266058 516986 266614
rect 517542 266058 517574 266614
rect 516954 230614 517574 266058
rect 516954 230058 516986 230614
rect 517542 230058 517574 230614
rect 516954 194614 517574 230058
rect 516954 194058 516986 194614
rect 517542 194058 517574 194614
rect 516954 158614 517574 194058
rect 516954 158058 516986 158614
rect 517542 158058 517574 158614
rect 516954 122614 517574 158058
rect 516954 122058 516986 122614
rect 517542 122058 517574 122614
rect 516954 86614 517574 122058
rect 516954 86058 516986 86614
rect 517542 86058 517574 86614
rect 516954 50614 517574 86058
rect 516954 50058 516986 50614
rect 517542 50058 517574 50614
rect 516954 14614 517574 50058
rect 516954 14058 516986 14614
rect 517542 14058 517574 14614
rect 516731 3500 516797 3501
rect 516731 3436 516732 3500
rect 516796 3436 516797 3500
rect 516731 3435 516797 3436
rect 514523 3228 514589 3229
rect 514523 3164 514524 3228
rect 514588 3164 514589 3228
rect 514523 3163 514589 3164
rect 514526 2821 514586 3163
rect 516734 2957 516794 3435
rect 516731 2956 516797 2957
rect 516731 2892 516732 2956
rect 516796 2892 516797 2956
rect 516731 2891 516797 2892
rect 514523 2820 514589 2821
rect 514523 2756 514524 2820
rect 514588 2756 514589 2820
rect 514523 2755 514589 2756
rect 513234 -2822 513266 -2266
rect 513822 -2822 513854 -2266
rect 513234 -7654 513854 -2822
rect 516954 -3226 517574 14058
rect 520674 708678 521294 711590
rect 520674 708122 520706 708678
rect 521262 708122 521294 708678
rect 520674 666334 521294 708122
rect 520674 665778 520706 666334
rect 521262 665778 521294 666334
rect 520674 630334 521294 665778
rect 520674 629778 520706 630334
rect 521262 629778 521294 630334
rect 520674 594334 521294 629778
rect 520674 593778 520706 594334
rect 521262 593778 521294 594334
rect 520674 558334 521294 593778
rect 520674 557778 520706 558334
rect 521262 557778 521294 558334
rect 520674 522334 521294 557778
rect 520674 521778 520706 522334
rect 521262 521778 521294 522334
rect 520674 486334 521294 521778
rect 520674 485778 520706 486334
rect 521262 485778 521294 486334
rect 520674 450334 521294 485778
rect 520674 449778 520706 450334
rect 521262 449778 521294 450334
rect 520674 414334 521294 449778
rect 520674 413778 520706 414334
rect 521262 413778 521294 414334
rect 520674 378334 521294 413778
rect 520674 377778 520706 378334
rect 521262 377778 521294 378334
rect 520674 342334 521294 377778
rect 520674 341778 520706 342334
rect 521262 341778 521294 342334
rect 520674 306334 521294 341778
rect 524394 709638 525014 711590
rect 524394 709082 524426 709638
rect 524982 709082 525014 709638
rect 524394 670054 525014 709082
rect 524394 669498 524426 670054
rect 524982 669498 525014 670054
rect 524394 634054 525014 669498
rect 524394 633498 524426 634054
rect 524982 633498 525014 634054
rect 524394 598054 525014 633498
rect 524394 597498 524426 598054
rect 524982 597498 525014 598054
rect 524394 562054 525014 597498
rect 524394 561498 524426 562054
rect 524982 561498 525014 562054
rect 524394 526054 525014 561498
rect 524394 525498 524426 526054
rect 524982 525498 525014 526054
rect 524394 490054 525014 525498
rect 524394 489498 524426 490054
rect 524982 489498 525014 490054
rect 524394 454054 525014 489498
rect 524394 453498 524426 454054
rect 524982 453498 525014 454054
rect 524394 418054 525014 453498
rect 524394 417498 524426 418054
rect 524982 417498 525014 418054
rect 524394 382054 525014 417498
rect 524394 381498 524426 382054
rect 524982 381498 525014 382054
rect 524394 346054 525014 381498
rect 524394 345498 524426 346054
rect 524982 345498 525014 346054
rect 523088 331174 523408 331206
rect 523088 330938 523130 331174
rect 523366 330938 523408 331174
rect 523088 330854 523408 330938
rect 523088 330618 523130 330854
rect 523366 330618 523408 330854
rect 523088 330586 523408 330618
rect 520674 305778 520706 306334
rect 521262 305778 521294 306334
rect 520674 270334 521294 305778
rect 524394 310054 525014 345498
rect 524394 309498 524426 310054
rect 524982 309498 525014 310054
rect 523088 295174 523408 295206
rect 523088 294938 523130 295174
rect 523366 294938 523408 295174
rect 523088 294854 523408 294938
rect 523088 294618 523130 294854
rect 523366 294618 523408 294854
rect 523088 294586 523408 294618
rect 520674 269778 520706 270334
rect 521262 269778 521294 270334
rect 520674 234334 521294 269778
rect 524394 274054 525014 309498
rect 524394 273498 524426 274054
rect 524982 273498 525014 274054
rect 523088 259174 523408 259206
rect 523088 258938 523130 259174
rect 523366 258938 523408 259174
rect 523088 258854 523408 258938
rect 523088 258618 523130 258854
rect 523366 258618 523408 258854
rect 523088 258586 523408 258618
rect 520674 233778 520706 234334
rect 521262 233778 521294 234334
rect 520674 198334 521294 233778
rect 524394 238054 525014 273498
rect 524394 237498 524426 238054
rect 524982 237498 525014 238054
rect 523088 223174 523408 223206
rect 523088 222938 523130 223174
rect 523366 222938 523408 223174
rect 523088 222854 523408 222938
rect 523088 222618 523130 222854
rect 523366 222618 523408 222854
rect 523088 222586 523408 222618
rect 520674 197778 520706 198334
rect 521262 197778 521294 198334
rect 520674 162334 521294 197778
rect 524394 202054 525014 237498
rect 524394 201498 524426 202054
rect 524982 201498 525014 202054
rect 523088 187174 523408 187206
rect 523088 186938 523130 187174
rect 523366 186938 523408 187174
rect 523088 186854 523408 186938
rect 523088 186618 523130 186854
rect 523366 186618 523408 186854
rect 523088 186586 523408 186618
rect 520674 161778 520706 162334
rect 521262 161778 521294 162334
rect 520674 126334 521294 161778
rect 524394 166054 525014 201498
rect 524394 165498 524426 166054
rect 524982 165498 525014 166054
rect 523088 151174 523408 151206
rect 523088 150938 523130 151174
rect 523366 150938 523408 151174
rect 523088 150854 523408 150938
rect 523088 150618 523130 150854
rect 523366 150618 523408 150854
rect 523088 150586 523408 150618
rect 520674 125778 520706 126334
rect 521262 125778 521294 126334
rect 520674 90334 521294 125778
rect 524394 130054 525014 165498
rect 524394 129498 524426 130054
rect 524982 129498 525014 130054
rect 523088 115174 523408 115206
rect 523088 114938 523130 115174
rect 523366 114938 523408 115174
rect 523088 114854 523408 114938
rect 523088 114618 523130 114854
rect 523366 114618 523408 114854
rect 523088 114586 523408 114618
rect 520674 89778 520706 90334
rect 521262 89778 521294 90334
rect 520674 54334 521294 89778
rect 524394 94054 525014 129498
rect 524394 93498 524426 94054
rect 524982 93498 525014 94054
rect 523088 79174 523408 79206
rect 523088 78938 523130 79174
rect 523366 78938 523408 79174
rect 523088 78854 523408 78938
rect 523088 78618 523130 78854
rect 523366 78618 523408 78854
rect 523088 78586 523408 78618
rect 520674 53778 520706 54334
rect 521262 53778 521294 54334
rect 520674 18334 521294 53778
rect 524394 58054 525014 93498
rect 524394 57498 524426 58054
rect 524982 57498 525014 58054
rect 523088 43174 523408 43206
rect 523088 42938 523130 43174
rect 523366 42938 523408 43174
rect 523088 42854 523408 42938
rect 523088 42618 523130 42854
rect 523366 42618 523408 42854
rect 523088 42586 523408 42618
rect 520674 17778 520706 18334
rect 521262 17778 521294 18334
rect 517835 3636 517901 3637
rect 517835 3572 517836 3636
rect 517900 3572 517901 3636
rect 517835 3571 517901 3572
rect 517838 3093 517898 3571
rect 517835 3092 517901 3093
rect 517835 3028 517836 3092
rect 517900 3028 517901 3092
rect 517835 3027 517901 3028
rect 516954 -3782 516986 -3226
rect 517542 -3782 517574 -3226
rect 516954 -7654 517574 -3782
rect 520674 -4186 521294 17778
rect 524394 22054 525014 57498
rect 524394 21498 524426 22054
rect 524982 21498 525014 22054
rect 523088 7174 523408 7206
rect 523088 6938 523130 7174
rect 523366 6938 523408 7174
rect 523088 6854 523408 6938
rect 523088 6618 523130 6854
rect 523366 6618 523408 6854
rect 523088 6586 523408 6618
rect 522987 3092 523053 3093
rect 522987 3028 522988 3092
rect 523052 3028 523053 3092
rect 522987 3027 523053 3028
rect 522990 2549 523050 3027
rect 522987 2548 523053 2549
rect 522987 2484 522988 2548
rect 523052 2484 523053 2548
rect 522987 2483 523053 2484
rect 520674 -4742 520706 -4186
rect 521262 -4742 521294 -4186
rect 520674 -7654 521294 -4742
rect 524394 -5146 525014 21498
rect 528114 710598 528734 711590
rect 528114 710042 528146 710598
rect 528702 710042 528734 710598
rect 528114 673774 528734 710042
rect 528114 673218 528146 673774
rect 528702 673218 528734 673774
rect 528114 637774 528734 673218
rect 528114 637218 528146 637774
rect 528702 637218 528734 637774
rect 528114 601774 528734 637218
rect 528114 601218 528146 601774
rect 528702 601218 528734 601774
rect 528114 565774 528734 601218
rect 528114 565218 528146 565774
rect 528702 565218 528734 565774
rect 528114 529774 528734 565218
rect 528114 529218 528146 529774
rect 528702 529218 528734 529774
rect 528114 493774 528734 529218
rect 528114 493218 528146 493774
rect 528702 493218 528734 493774
rect 528114 457774 528734 493218
rect 528114 457218 528146 457774
rect 528702 457218 528734 457774
rect 528114 421774 528734 457218
rect 528114 421218 528146 421774
rect 528702 421218 528734 421774
rect 528114 385774 528734 421218
rect 528114 385218 528146 385774
rect 528702 385218 528734 385774
rect 528114 349774 528734 385218
rect 528114 349218 528146 349774
rect 528702 349218 528734 349774
rect 528114 313774 528734 349218
rect 528114 313218 528146 313774
rect 528702 313218 528734 313774
rect 528114 277774 528734 313218
rect 528114 277218 528146 277774
rect 528702 277218 528734 277774
rect 528114 241774 528734 277218
rect 528114 241218 528146 241774
rect 528702 241218 528734 241774
rect 528114 205774 528734 241218
rect 528114 205218 528146 205774
rect 528702 205218 528734 205774
rect 528114 169774 528734 205218
rect 528114 169218 528146 169774
rect 528702 169218 528734 169774
rect 528114 133774 528734 169218
rect 528114 133218 528146 133774
rect 528702 133218 528734 133774
rect 528114 97774 528734 133218
rect 528114 97218 528146 97774
rect 528702 97218 528734 97774
rect 528114 61774 528734 97218
rect 528114 61218 528146 61774
rect 528702 61218 528734 61774
rect 528114 25774 528734 61218
rect 528114 25218 528146 25774
rect 528702 25218 528734 25774
rect 526299 3636 526365 3637
rect 526299 3572 526300 3636
rect 526364 3572 526365 3636
rect 526299 3571 526365 3572
rect 526302 2957 526362 3571
rect 526483 3092 526549 3093
rect 526483 3028 526484 3092
rect 526548 3028 526549 3092
rect 526483 3027 526549 3028
rect 527587 3092 527653 3093
rect 527587 3028 527588 3092
rect 527652 3028 527653 3092
rect 527587 3027 527653 3028
rect 526299 2956 526365 2957
rect 526299 2892 526300 2956
rect 526364 2892 526365 2956
rect 526299 2891 526365 2892
rect 526486 2685 526546 3027
rect 527590 2685 527650 3027
rect 526483 2684 526549 2685
rect 526483 2620 526484 2684
rect 526548 2620 526549 2684
rect 526483 2619 526549 2620
rect 527587 2684 527653 2685
rect 527587 2620 527588 2684
rect 527652 2620 527653 2684
rect 527587 2619 527653 2620
rect 524394 -5702 524426 -5146
rect 524982 -5702 525014 -5146
rect 524394 -7654 525014 -5702
rect 528114 -6106 528734 25218
rect 531834 711558 532454 711590
rect 531834 711002 531866 711558
rect 532422 711002 532454 711558
rect 531834 677494 532454 711002
rect 531834 676938 531866 677494
rect 532422 676938 532454 677494
rect 531834 641494 532454 676938
rect 531834 640938 531866 641494
rect 532422 640938 532454 641494
rect 531834 605494 532454 640938
rect 531834 604938 531866 605494
rect 532422 604938 532454 605494
rect 531834 569494 532454 604938
rect 531834 568938 531866 569494
rect 532422 568938 532454 569494
rect 531834 533494 532454 568938
rect 531834 532938 531866 533494
rect 532422 532938 532454 533494
rect 531834 497494 532454 532938
rect 531834 496938 531866 497494
rect 532422 496938 532454 497494
rect 531834 461494 532454 496938
rect 531834 460938 531866 461494
rect 532422 460938 532454 461494
rect 531834 425494 532454 460938
rect 531834 424938 531866 425494
rect 532422 424938 532454 425494
rect 531834 389494 532454 424938
rect 531834 388938 531866 389494
rect 532422 388938 532454 389494
rect 531834 353494 532454 388938
rect 531834 352938 531866 353494
rect 532422 352938 532454 353494
rect 531834 317494 532454 352938
rect 541794 704838 542414 711590
rect 541794 704282 541826 704838
rect 542382 704282 542414 704838
rect 541794 687454 542414 704282
rect 541794 686898 541826 687454
rect 542382 686898 542414 687454
rect 541794 651454 542414 686898
rect 541794 650898 541826 651454
rect 542382 650898 542414 651454
rect 541794 615454 542414 650898
rect 541794 614898 541826 615454
rect 542382 614898 542414 615454
rect 541794 579454 542414 614898
rect 541794 578898 541826 579454
rect 542382 578898 542414 579454
rect 541794 543454 542414 578898
rect 541794 542898 541826 543454
rect 542382 542898 542414 543454
rect 541794 507454 542414 542898
rect 541794 506898 541826 507454
rect 542382 506898 542414 507454
rect 541794 471454 542414 506898
rect 541794 470898 541826 471454
rect 542382 470898 542414 471454
rect 541794 435454 542414 470898
rect 541794 434898 541826 435454
rect 542382 434898 542414 435454
rect 541794 399454 542414 434898
rect 541794 398898 541826 399454
rect 542382 398898 542414 399454
rect 541794 363454 542414 398898
rect 541794 362898 541826 363454
rect 542382 362898 542414 363454
rect 538448 327454 538768 327486
rect 538448 327218 538490 327454
rect 538726 327218 538768 327454
rect 538448 327134 538768 327218
rect 538448 326898 538490 327134
rect 538726 326898 538768 327134
rect 538448 326866 538768 326898
rect 541794 327454 542414 362898
rect 541794 326898 541826 327454
rect 542382 326898 542414 327454
rect 531834 316938 531866 317494
rect 532422 316938 532454 317494
rect 531834 281494 532454 316938
rect 538448 291454 538768 291486
rect 538448 291218 538490 291454
rect 538726 291218 538768 291454
rect 538448 291134 538768 291218
rect 538448 290898 538490 291134
rect 538726 290898 538768 291134
rect 538448 290866 538768 290898
rect 541794 291454 542414 326898
rect 541794 290898 541826 291454
rect 542382 290898 542414 291454
rect 531834 280938 531866 281494
rect 532422 280938 532454 281494
rect 531834 245494 532454 280938
rect 538448 255454 538768 255486
rect 538448 255218 538490 255454
rect 538726 255218 538768 255454
rect 538448 255134 538768 255218
rect 538448 254898 538490 255134
rect 538726 254898 538768 255134
rect 538448 254866 538768 254898
rect 541794 255454 542414 290898
rect 541794 254898 541826 255454
rect 542382 254898 542414 255454
rect 531834 244938 531866 245494
rect 532422 244938 532454 245494
rect 531834 209494 532454 244938
rect 538448 219454 538768 219486
rect 538448 219218 538490 219454
rect 538726 219218 538768 219454
rect 538448 219134 538768 219218
rect 538448 218898 538490 219134
rect 538726 218898 538768 219134
rect 538448 218866 538768 218898
rect 541794 219454 542414 254898
rect 541794 218898 541826 219454
rect 542382 218898 542414 219454
rect 531834 208938 531866 209494
rect 532422 208938 532454 209494
rect 531834 173494 532454 208938
rect 538448 183454 538768 183486
rect 538448 183218 538490 183454
rect 538726 183218 538768 183454
rect 538448 183134 538768 183218
rect 538448 182898 538490 183134
rect 538726 182898 538768 183134
rect 538448 182866 538768 182898
rect 541794 183454 542414 218898
rect 541794 182898 541826 183454
rect 542382 182898 542414 183454
rect 531834 172938 531866 173494
rect 532422 172938 532454 173494
rect 531834 137494 532454 172938
rect 538448 147454 538768 147486
rect 538448 147218 538490 147454
rect 538726 147218 538768 147454
rect 538448 147134 538768 147218
rect 538448 146898 538490 147134
rect 538726 146898 538768 147134
rect 538448 146866 538768 146898
rect 541794 147454 542414 182898
rect 541794 146898 541826 147454
rect 542382 146898 542414 147454
rect 531834 136938 531866 137494
rect 532422 136938 532454 137494
rect 531834 101494 532454 136938
rect 538448 111454 538768 111486
rect 538448 111218 538490 111454
rect 538726 111218 538768 111454
rect 538448 111134 538768 111218
rect 538448 110898 538490 111134
rect 538726 110898 538768 111134
rect 538448 110866 538768 110898
rect 541794 111454 542414 146898
rect 541794 110898 541826 111454
rect 542382 110898 542414 111454
rect 531834 100938 531866 101494
rect 532422 100938 532454 101494
rect 531834 65494 532454 100938
rect 538448 75454 538768 75486
rect 538448 75218 538490 75454
rect 538726 75218 538768 75454
rect 538448 75134 538768 75218
rect 538448 74898 538490 75134
rect 538726 74898 538768 75134
rect 538448 74866 538768 74898
rect 541794 75454 542414 110898
rect 541794 74898 541826 75454
rect 542382 74898 542414 75454
rect 531834 64938 531866 65494
rect 532422 64938 532454 65494
rect 531834 29494 532454 64938
rect 538448 39454 538768 39486
rect 538448 39218 538490 39454
rect 538726 39218 538768 39454
rect 538448 39134 538768 39218
rect 538448 38898 538490 39134
rect 538726 38898 538768 39134
rect 538448 38866 538768 38898
rect 541794 39454 542414 74898
rect 541794 38898 541826 39454
rect 542382 38898 542414 39454
rect 531834 28938 531866 29494
rect 532422 28938 532454 29494
rect 529979 3228 530045 3229
rect 529979 3164 529980 3228
rect 530044 3164 530045 3228
rect 529979 3163 530045 3164
rect 529982 2685 530042 3163
rect 529979 2684 530045 2685
rect 529979 2620 529980 2684
rect 530044 2620 530045 2684
rect 529979 2619 530045 2620
rect 528114 -6662 528146 -6106
rect 528702 -6662 528734 -6106
rect 528114 -7654 528734 -6662
rect 531834 -7066 532454 28938
rect 533475 3772 533541 3773
rect 533475 3708 533476 3772
rect 533540 3708 533541 3772
rect 533475 3707 533541 3708
rect 533478 2957 533538 3707
rect 541794 3454 542414 38898
rect 545514 705798 546134 711590
rect 545514 705242 545546 705798
rect 546102 705242 546134 705798
rect 545514 691174 546134 705242
rect 545514 690618 545546 691174
rect 546102 690618 546134 691174
rect 545514 655174 546134 690618
rect 545514 654618 545546 655174
rect 546102 654618 546134 655174
rect 545514 619174 546134 654618
rect 545514 618618 545546 619174
rect 546102 618618 546134 619174
rect 545514 583174 546134 618618
rect 545514 582618 545546 583174
rect 546102 582618 546134 583174
rect 545514 547174 546134 582618
rect 545514 546618 545546 547174
rect 546102 546618 546134 547174
rect 545514 511174 546134 546618
rect 545514 510618 545546 511174
rect 546102 510618 546134 511174
rect 545514 475174 546134 510618
rect 545514 474618 545546 475174
rect 546102 474618 546134 475174
rect 545514 439174 546134 474618
rect 545514 438618 545546 439174
rect 546102 438618 546134 439174
rect 545514 403174 546134 438618
rect 545514 402618 545546 403174
rect 546102 402618 546134 403174
rect 545514 367174 546134 402618
rect 545514 366618 545546 367174
rect 546102 366618 546134 367174
rect 545514 331174 546134 366618
rect 545514 330618 545546 331174
rect 546102 330618 546134 331174
rect 545514 295174 546134 330618
rect 545514 294618 545546 295174
rect 546102 294618 546134 295174
rect 545514 259174 546134 294618
rect 545514 258618 545546 259174
rect 546102 258618 546134 259174
rect 545514 223174 546134 258618
rect 545514 222618 545546 223174
rect 546102 222618 546134 223174
rect 545514 187174 546134 222618
rect 545514 186618 545546 187174
rect 546102 186618 546134 187174
rect 545514 151174 546134 186618
rect 545514 150618 545546 151174
rect 546102 150618 546134 151174
rect 545514 115174 546134 150618
rect 545514 114618 545546 115174
rect 546102 114618 546134 115174
rect 545514 79174 546134 114618
rect 545514 78618 545546 79174
rect 546102 78618 546134 79174
rect 545514 43174 546134 78618
rect 545514 42618 545546 43174
rect 546102 42618 546134 43174
rect 545514 7174 546134 42618
rect 545514 6618 545546 7174
rect 546102 6618 546134 7174
rect 545251 3636 545317 3637
rect 545251 3572 545252 3636
rect 545316 3572 545317 3636
rect 545251 3571 545317 3572
rect 533475 2956 533541 2957
rect 533475 2892 533476 2956
rect 533540 2892 533541 2956
rect 533475 2891 533541 2892
rect 541794 2898 541826 3454
rect 542382 2898 542414 3454
rect 533291 2820 533357 2821
rect 533291 2756 533292 2820
rect 533356 2756 533357 2820
rect 533291 2755 533357 2756
rect 533294 2685 533354 2755
rect 533291 2684 533357 2685
rect 533291 2620 533292 2684
rect 533356 2620 533357 2684
rect 533291 2619 533357 2620
rect 531834 -7622 531866 -7066
rect 532422 -7622 532454 -7066
rect 531834 -7654 532454 -7622
rect 541794 -346 542414 2898
rect 545254 2549 545314 3571
rect 545251 2548 545317 2549
rect 545251 2484 545252 2548
rect 545316 2484 545317 2548
rect 545251 2483 545317 2484
rect 541794 -902 541826 -346
rect 542382 -902 542414 -346
rect 541794 -7654 542414 -902
rect 545514 -1306 546134 6618
rect 549234 706758 549854 711590
rect 549234 706202 549266 706758
rect 549822 706202 549854 706758
rect 549234 694894 549854 706202
rect 549234 694338 549266 694894
rect 549822 694338 549854 694894
rect 549234 658894 549854 694338
rect 549234 658338 549266 658894
rect 549822 658338 549854 658894
rect 549234 622894 549854 658338
rect 549234 622338 549266 622894
rect 549822 622338 549854 622894
rect 549234 586894 549854 622338
rect 549234 586338 549266 586894
rect 549822 586338 549854 586894
rect 549234 550894 549854 586338
rect 549234 550338 549266 550894
rect 549822 550338 549854 550894
rect 549234 514894 549854 550338
rect 549234 514338 549266 514894
rect 549822 514338 549854 514894
rect 549234 478894 549854 514338
rect 549234 478338 549266 478894
rect 549822 478338 549854 478894
rect 549234 442894 549854 478338
rect 549234 442338 549266 442894
rect 549822 442338 549854 442894
rect 549234 406894 549854 442338
rect 549234 406338 549266 406894
rect 549822 406338 549854 406894
rect 549234 370894 549854 406338
rect 549234 370338 549266 370894
rect 549822 370338 549854 370894
rect 549234 334894 549854 370338
rect 549234 334338 549266 334894
rect 549822 334338 549854 334894
rect 549234 298894 549854 334338
rect 549234 298338 549266 298894
rect 549822 298338 549854 298894
rect 549234 262894 549854 298338
rect 549234 262338 549266 262894
rect 549822 262338 549854 262894
rect 549234 226894 549854 262338
rect 549234 226338 549266 226894
rect 549822 226338 549854 226894
rect 549234 190894 549854 226338
rect 549234 190338 549266 190894
rect 549822 190338 549854 190894
rect 549234 154894 549854 190338
rect 549234 154338 549266 154894
rect 549822 154338 549854 154894
rect 549234 118894 549854 154338
rect 549234 118338 549266 118894
rect 549822 118338 549854 118894
rect 549234 82894 549854 118338
rect 549234 82338 549266 82894
rect 549822 82338 549854 82894
rect 549234 46894 549854 82338
rect 549234 46338 549266 46894
rect 549822 46338 549854 46894
rect 549234 10894 549854 46338
rect 549234 10338 549266 10894
rect 549822 10338 549854 10894
rect 547643 3500 547709 3501
rect 547643 3436 547644 3500
rect 547708 3436 547709 3500
rect 547643 3435 547709 3436
rect 547646 2549 547706 3435
rect 547643 2548 547709 2549
rect 547643 2484 547644 2548
rect 547708 2484 547709 2548
rect 547643 2483 547709 2484
rect 545514 -1862 545546 -1306
rect 546102 -1862 546134 -1306
rect 545514 -7654 546134 -1862
rect 549234 -2266 549854 10338
rect 552954 707718 553574 711590
rect 552954 707162 552986 707718
rect 553542 707162 553574 707718
rect 552954 698614 553574 707162
rect 552954 698058 552986 698614
rect 553542 698058 553574 698614
rect 552954 662614 553574 698058
rect 552954 662058 552986 662614
rect 553542 662058 553574 662614
rect 552954 626614 553574 662058
rect 552954 626058 552986 626614
rect 553542 626058 553574 626614
rect 552954 590614 553574 626058
rect 552954 590058 552986 590614
rect 553542 590058 553574 590614
rect 552954 554614 553574 590058
rect 552954 554058 552986 554614
rect 553542 554058 553574 554614
rect 552954 518614 553574 554058
rect 552954 518058 552986 518614
rect 553542 518058 553574 518614
rect 552954 482614 553574 518058
rect 552954 482058 552986 482614
rect 553542 482058 553574 482614
rect 552954 446614 553574 482058
rect 552954 446058 552986 446614
rect 553542 446058 553574 446614
rect 552954 410614 553574 446058
rect 552954 410058 552986 410614
rect 553542 410058 553574 410614
rect 552954 374614 553574 410058
rect 552954 374058 552986 374614
rect 553542 374058 553574 374614
rect 552954 338614 553574 374058
rect 552954 338058 552986 338614
rect 553542 338058 553574 338614
rect 552954 302614 553574 338058
rect 556674 708678 557294 711590
rect 556674 708122 556706 708678
rect 557262 708122 557294 708678
rect 556674 666334 557294 708122
rect 556674 665778 556706 666334
rect 557262 665778 557294 666334
rect 556674 630334 557294 665778
rect 556674 629778 556706 630334
rect 557262 629778 557294 630334
rect 556674 594334 557294 629778
rect 556674 593778 556706 594334
rect 557262 593778 557294 594334
rect 556674 558334 557294 593778
rect 556674 557778 556706 558334
rect 557262 557778 557294 558334
rect 556674 522334 557294 557778
rect 556674 521778 556706 522334
rect 557262 521778 557294 522334
rect 556674 486334 557294 521778
rect 556674 485778 556706 486334
rect 557262 485778 557294 486334
rect 556674 450334 557294 485778
rect 556674 449778 556706 450334
rect 557262 449778 557294 450334
rect 556674 414334 557294 449778
rect 556674 413778 556706 414334
rect 557262 413778 557294 414334
rect 556674 378334 557294 413778
rect 556674 377778 556706 378334
rect 557262 377778 557294 378334
rect 556674 342334 557294 377778
rect 556674 341778 556706 342334
rect 557262 341778 557294 342334
rect 553808 331174 554128 331206
rect 553808 330938 553850 331174
rect 554086 330938 554128 331174
rect 553808 330854 554128 330938
rect 553808 330618 553850 330854
rect 554086 330618 554128 330854
rect 553808 330586 554128 330618
rect 552954 302058 552986 302614
rect 553542 302058 553574 302614
rect 552954 266614 553574 302058
rect 556674 306334 557294 341778
rect 556674 305778 556706 306334
rect 557262 305778 557294 306334
rect 553808 295174 554128 295206
rect 553808 294938 553850 295174
rect 554086 294938 554128 295174
rect 553808 294854 554128 294938
rect 553808 294618 553850 294854
rect 554086 294618 554128 294854
rect 553808 294586 554128 294618
rect 552954 266058 552986 266614
rect 553542 266058 553574 266614
rect 552954 230614 553574 266058
rect 556674 270334 557294 305778
rect 556674 269778 556706 270334
rect 557262 269778 557294 270334
rect 553808 259174 554128 259206
rect 553808 258938 553850 259174
rect 554086 258938 554128 259174
rect 553808 258854 554128 258938
rect 553808 258618 553850 258854
rect 554086 258618 554128 258854
rect 553808 258586 554128 258618
rect 552954 230058 552986 230614
rect 553542 230058 553574 230614
rect 552954 194614 553574 230058
rect 556674 234334 557294 269778
rect 556674 233778 556706 234334
rect 557262 233778 557294 234334
rect 553808 223174 554128 223206
rect 553808 222938 553850 223174
rect 554086 222938 554128 223174
rect 553808 222854 554128 222938
rect 553808 222618 553850 222854
rect 554086 222618 554128 222854
rect 553808 222586 554128 222618
rect 552954 194058 552986 194614
rect 553542 194058 553574 194614
rect 552954 158614 553574 194058
rect 556674 198334 557294 233778
rect 556674 197778 556706 198334
rect 557262 197778 557294 198334
rect 553808 187174 554128 187206
rect 553808 186938 553850 187174
rect 554086 186938 554128 187174
rect 553808 186854 554128 186938
rect 553808 186618 553850 186854
rect 554086 186618 554128 186854
rect 553808 186586 554128 186618
rect 552954 158058 552986 158614
rect 553542 158058 553574 158614
rect 552954 122614 553574 158058
rect 556674 162334 557294 197778
rect 556674 161778 556706 162334
rect 557262 161778 557294 162334
rect 553808 151174 554128 151206
rect 553808 150938 553850 151174
rect 554086 150938 554128 151174
rect 553808 150854 554128 150938
rect 553808 150618 553850 150854
rect 554086 150618 554128 150854
rect 553808 150586 554128 150618
rect 552954 122058 552986 122614
rect 553542 122058 553574 122614
rect 552954 86614 553574 122058
rect 556674 126334 557294 161778
rect 556674 125778 556706 126334
rect 557262 125778 557294 126334
rect 553808 115174 554128 115206
rect 553808 114938 553850 115174
rect 554086 114938 554128 115174
rect 553808 114854 554128 114938
rect 553808 114618 553850 114854
rect 554086 114618 554128 114854
rect 553808 114586 554128 114618
rect 552954 86058 552986 86614
rect 553542 86058 553574 86614
rect 552954 50614 553574 86058
rect 556674 90334 557294 125778
rect 556674 89778 556706 90334
rect 557262 89778 557294 90334
rect 553808 79174 554128 79206
rect 553808 78938 553850 79174
rect 554086 78938 554128 79174
rect 553808 78854 554128 78938
rect 553808 78618 553850 78854
rect 554086 78618 554128 78854
rect 553808 78586 554128 78618
rect 552954 50058 552986 50614
rect 553542 50058 553574 50614
rect 552954 14614 553574 50058
rect 556674 54334 557294 89778
rect 556674 53778 556706 54334
rect 557262 53778 557294 54334
rect 553808 43174 554128 43206
rect 553808 42938 553850 43174
rect 554086 42938 554128 43174
rect 553808 42854 554128 42938
rect 553808 42618 553850 42854
rect 554086 42618 554128 42854
rect 553808 42586 554128 42618
rect 552954 14058 552986 14614
rect 553542 14058 553574 14614
rect 552427 3364 552493 3365
rect 552427 3300 552428 3364
rect 552492 3300 552493 3364
rect 552427 3299 552493 3300
rect 552430 2685 552490 3299
rect 552427 2684 552493 2685
rect 552427 2620 552428 2684
rect 552492 2620 552493 2684
rect 552427 2619 552493 2620
rect 549234 -2822 549266 -2266
rect 549822 -2822 549854 -2266
rect 549234 -7654 549854 -2822
rect 552954 -3226 553574 14058
rect 556674 18334 557294 53778
rect 556674 17778 556706 18334
rect 557262 17778 557294 18334
rect 553808 7174 554128 7206
rect 553808 6938 553850 7174
rect 554086 6938 554128 7174
rect 553808 6854 554128 6938
rect 553808 6618 553850 6854
rect 554086 6618 554128 6854
rect 553808 6586 554128 6618
rect 552954 -3782 552986 -3226
rect 553542 -3782 553574 -3226
rect 552954 -7654 553574 -3782
rect 556674 -4186 557294 17778
rect 560394 709638 561014 711590
rect 560394 709082 560426 709638
rect 560982 709082 561014 709638
rect 560394 670054 561014 709082
rect 560394 669498 560426 670054
rect 560982 669498 561014 670054
rect 560394 634054 561014 669498
rect 560394 633498 560426 634054
rect 560982 633498 561014 634054
rect 560394 598054 561014 633498
rect 560394 597498 560426 598054
rect 560982 597498 561014 598054
rect 560394 562054 561014 597498
rect 560394 561498 560426 562054
rect 560982 561498 561014 562054
rect 560394 526054 561014 561498
rect 560394 525498 560426 526054
rect 560982 525498 561014 526054
rect 560394 490054 561014 525498
rect 560394 489498 560426 490054
rect 560982 489498 561014 490054
rect 560394 454054 561014 489498
rect 560394 453498 560426 454054
rect 560982 453498 561014 454054
rect 560394 418054 561014 453498
rect 560394 417498 560426 418054
rect 560982 417498 561014 418054
rect 560394 382054 561014 417498
rect 560394 381498 560426 382054
rect 560982 381498 561014 382054
rect 560394 346054 561014 381498
rect 560394 345498 560426 346054
rect 560982 345498 561014 346054
rect 560394 310054 561014 345498
rect 560394 309498 560426 310054
rect 560982 309498 561014 310054
rect 560394 274054 561014 309498
rect 560394 273498 560426 274054
rect 560982 273498 561014 274054
rect 560394 238054 561014 273498
rect 560394 237498 560426 238054
rect 560982 237498 561014 238054
rect 560394 202054 561014 237498
rect 560394 201498 560426 202054
rect 560982 201498 561014 202054
rect 560394 166054 561014 201498
rect 560394 165498 560426 166054
rect 560982 165498 561014 166054
rect 560394 130054 561014 165498
rect 560394 129498 560426 130054
rect 560982 129498 561014 130054
rect 560394 94054 561014 129498
rect 560394 93498 560426 94054
rect 560982 93498 561014 94054
rect 560394 58054 561014 93498
rect 560394 57498 560426 58054
rect 560982 57498 561014 58054
rect 560394 22054 561014 57498
rect 560394 21498 560426 22054
rect 560982 21498 561014 22054
rect 558499 3908 558565 3909
rect 558499 3844 558500 3908
rect 558564 3844 558565 3908
rect 558499 3843 558565 3844
rect 558502 2821 558562 3843
rect 558499 2820 558565 2821
rect 558499 2756 558500 2820
rect 558564 2756 558565 2820
rect 558499 2755 558565 2756
rect 556674 -4742 556706 -4186
rect 557262 -4742 557294 -4186
rect 556674 -7654 557294 -4742
rect 560394 -5146 561014 21498
rect 560394 -5702 560426 -5146
rect 560982 -5702 561014 -5146
rect 560394 -7654 561014 -5702
rect 564114 710598 564734 711590
rect 564114 710042 564146 710598
rect 564702 710042 564734 710598
rect 564114 673774 564734 710042
rect 564114 673218 564146 673774
rect 564702 673218 564734 673774
rect 564114 637774 564734 673218
rect 564114 637218 564146 637774
rect 564702 637218 564734 637774
rect 564114 601774 564734 637218
rect 564114 601218 564146 601774
rect 564702 601218 564734 601774
rect 564114 565774 564734 601218
rect 564114 565218 564146 565774
rect 564702 565218 564734 565774
rect 564114 529774 564734 565218
rect 564114 529218 564146 529774
rect 564702 529218 564734 529774
rect 564114 493774 564734 529218
rect 564114 493218 564146 493774
rect 564702 493218 564734 493774
rect 564114 457774 564734 493218
rect 564114 457218 564146 457774
rect 564702 457218 564734 457774
rect 564114 421774 564734 457218
rect 564114 421218 564146 421774
rect 564702 421218 564734 421774
rect 564114 385774 564734 421218
rect 564114 385218 564146 385774
rect 564702 385218 564734 385774
rect 564114 349774 564734 385218
rect 564114 349218 564146 349774
rect 564702 349218 564734 349774
rect 564114 313774 564734 349218
rect 564114 313218 564146 313774
rect 564702 313218 564734 313774
rect 564114 277774 564734 313218
rect 564114 277218 564146 277774
rect 564702 277218 564734 277774
rect 564114 241774 564734 277218
rect 564114 241218 564146 241774
rect 564702 241218 564734 241774
rect 564114 205774 564734 241218
rect 564114 205218 564146 205774
rect 564702 205218 564734 205774
rect 564114 169774 564734 205218
rect 564114 169218 564146 169774
rect 564702 169218 564734 169774
rect 564114 133774 564734 169218
rect 564114 133218 564146 133774
rect 564702 133218 564734 133774
rect 564114 97774 564734 133218
rect 564114 97218 564146 97774
rect 564702 97218 564734 97774
rect 564114 61774 564734 97218
rect 564114 61218 564146 61774
rect 564702 61218 564734 61774
rect 564114 25774 564734 61218
rect 564114 25218 564146 25774
rect 564702 25218 564734 25774
rect 564114 -6106 564734 25218
rect 564114 -6662 564146 -6106
rect 564702 -6662 564734 -6106
rect 564114 -7654 564734 -6662
rect 567834 711558 568454 711590
rect 567834 711002 567866 711558
rect 568422 711002 568454 711558
rect 567834 677494 568454 711002
rect 567834 676938 567866 677494
rect 568422 676938 568454 677494
rect 567834 641494 568454 676938
rect 567834 640938 567866 641494
rect 568422 640938 568454 641494
rect 567834 605494 568454 640938
rect 567834 604938 567866 605494
rect 568422 604938 568454 605494
rect 567834 569494 568454 604938
rect 567834 568938 567866 569494
rect 568422 568938 568454 569494
rect 567834 533494 568454 568938
rect 567834 532938 567866 533494
rect 568422 532938 568454 533494
rect 567834 497494 568454 532938
rect 567834 496938 567866 497494
rect 568422 496938 568454 497494
rect 567834 461494 568454 496938
rect 567834 460938 567866 461494
rect 568422 460938 568454 461494
rect 567834 425494 568454 460938
rect 567834 424938 567866 425494
rect 568422 424938 568454 425494
rect 567834 389494 568454 424938
rect 567834 388938 567866 389494
rect 568422 388938 568454 389494
rect 567834 353494 568454 388938
rect 567834 352938 567866 353494
rect 568422 352938 568454 353494
rect 567834 317494 568454 352938
rect 577794 704838 578414 711590
rect 577794 704282 577826 704838
rect 578382 704282 578414 704838
rect 577794 687454 578414 704282
rect 577794 686898 577826 687454
rect 578382 686898 578414 687454
rect 577794 651454 578414 686898
rect 577794 650898 577826 651454
rect 578382 650898 578414 651454
rect 577794 615454 578414 650898
rect 577794 614898 577826 615454
rect 578382 614898 578414 615454
rect 577794 579454 578414 614898
rect 577794 578898 577826 579454
rect 578382 578898 578414 579454
rect 577794 543454 578414 578898
rect 577794 542898 577826 543454
rect 578382 542898 578414 543454
rect 577794 507454 578414 542898
rect 577794 506898 577826 507454
rect 578382 506898 578414 507454
rect 577794 471454 578414 506898
rect 577794 470898 577826 471454
rect 578382 470898 578414 471454
rect 577794 435454 578414 470898
rect 577794 434898 577826 435454
rect 578382 434898 578414 435454
rect 577794 399454 578414 434898
rect 577794 398898 577826 399454
rect 578382 398898 578414 399454
rect 577794 363454 578414 398898
rect 577794 362898 577826 363454
rect 578382 362898 578414 363454
rect 574691 344724 574757 344725
rect 574691 344660 574692 344724
rect 574756 344660 574757 344724
rect 574691 344659 574757 344660
rect 569168 327454 569488 327486
rect 569168 327218 569210 327454
rect 569446 327218 569488 327454
rect 569168 327134 569488 327218
rect 569168 326898 569210 327134
rect 569446 326898 569488 327134
rect 569168 326866 569488 326898
rect 574694 325277 574754 344659
rect 574875 330308 574941 330309
rect 574875 330244 574876 330308
rect 574940 330244 574941 330308
rect 574875 330243 574941 330244
rect 574691 325276 574757 325277
rect 574691 325212 574692 325276
rect 574756 325212 574757 325276
rect 574691 325211 574757 325212
rect 567834 316938 567866 317494
rect 568422 316938 568454 317494
rect 567834 281494 568454 316938
rect 574878 312085 574938 330243
rect 577794 327454 578414 362898
rect 577794 326898 577826 327454
rect 578382 326898 578414 327454
rect 575059 315892 575125 315893
rect 575059 315828 575060 315892
rect 575124 315828 575125 315892
rect 575059 315827 575125 315828
rect 574875 312084 574941 312085
rect 574875 312020 574876 312084
rect 574940 312020 574941 312084
rect 574875 312019 574941 312020
rect 574691 301476 574757 301477
rect 574691 301412 574692 301476
rect 574756 301412 574757 301476
rect 574691 301411 574757 301412
rect 569168 291454 569488 291486
rect 569168 291218 569210 291454
rect 569446 291218 569488 291454
rect 569168 291134 569488 291218
rect 569168 290898 569210 291134
rect 569446 290898 569488 291134
rect 569168 290866 569488 290898
rect 567834 280938 567866 281494
rect 568422 280938 568454 281494
rect 567834 245494 568454 280938
rect 574694 272237 574754 301411
rect 575062 298757 575122 315827
rect 575059 298756 575125 298757
rect 575059 298692 575060 298756
rect 575124 298692 575125 298756
rect 575059 298691 575125 298692
rect 577794 291454 578414 326898
rect 577794 290898 577826 291454
rect 578382 290898 578414 291454
rect 575059 287060 575125 287061
rect 575059 286996 575060 287060
rect 575124 286996 575125 287060
rect 575059 286995 575125 286996
rect 574875 272644 574941 272645
rect 574875 272580 574876 272644
rect 574940 272580 574941 272644
rect 574875 272579 574941 272580
rect 574691 272236 574757 272237
rect 574691 272172 574692 272236
rect 574756 272172 574757 272236
rect 574691 272171 574757 272172
rect 574691 258228 574757 258229
rect 574691 258164 574692 258228
rect 574756 258164 574757 258228
rect 574691 258163 574757 258164
rect 569168 255454 569488 255486
rect 569168 255218 569210 255454
rect 569446 255218 569488 255454
rect 569168 255134 569488 255218
rect 569168 254898 569210 255134
rect 569446 254898 569488 255134
rect 569168 254866 569488 254898
rect 567834 244938 567866 245494
rect 568422 244938 568454 245494
rect 567834 209494 568454 244938
rect 574694 232389 574754 258163
rect 574878 245581 574938 272579
rect 575062 258909 575122 286995
rect 575059 258908 575125 258909
rect 575059 258844 575060 258908
rect 575124 258844 575125 258908
rect 575059 258843 575125 258844
rect 577794 255454 578414 290898
rect 577794 254898 577826 255454
rect 578382 254898 578414 255454
rect 574875 245580 574941 245581
rect 574875 245516 574876 245580
rect 574940 245516 574941 245580
rect 574875 245515 574941 245516
rect 574875 243812 574941 243813
rect 574875 243748 574876 243812
rect 574940 243748 574941 243812
rect 574875 243747 574941 243748
rect 574691 232388 574757 232389
rect 574691 232324 574692 232388
rect 574756 232324 574757 232388
rect 574691 232323 574757 232324
rect 574691 229396 574757 229397
rect 574691 229332 574692 229396
rect 574756 229332 574757 229396
rect 574691 229331 574757 229332
rect 569168 219454 569488 219486
rect 569168 219218 569210 219454
rect 569446 219218 569488 219454
rect 569168 219134 569488 219218
rect 569168 218898 569210 219134
rect 569446 218898 569488 219134
rect 569168 218866 569488 218898
rect 567834 208938 567866 209494
rect 568422 208938 568454 209494
rect 567834 173494 568454 208938
rect 574694 205733 574754 229331
rect 574878 219061 574938 243747
rect 577794 219454 578414 254898
rect 574875 219060 574941 219061
rect 574875 218996 574876 219060
rect 574940 218996 574941 219060
rect 574875 218995 574941 218996
rect 577794 218898 577826 219454
rect 578382 218898 578414 219454
rect 574875 214980 574941 214981
rect 574875 214916 574876 214980
rect 574940 214916 574941 214980
rect 574875 214915 574941 214916
rect 574691 205732 574757 205733
rect 574691 205668 574692 205732
rect 574756 205668 574757 205732
rect 574691 205667 574757 205668
rect 574691 200564 574757 200565
rect 574691 200500 574692 200564
rect 574756 200500 574757 200564
rect 574691 200499 574757 200500
rect 569168 183454 569488 183486
rect 569168 183218 569210 183454
rect 569446 183218 569488 183454
rect 569168 183134 569488 183218
rect 569168 182898 569210 183134
rect 569446 182898 569488 183134
rect 569168 182866 569488 182898
rect 574694 179213 574754 200499
rect 574878 192541 574938 214915
rect 574875 192540 574941 192541
rect 574875 192476 574876 192540
rect 574940 192476 574941 192540
rect 574875 192475 574941 192476
rect 574875 186148 574941 186149
rect 574875 186084 574876 186148
rect 574940 186084 574941 186148
rect 574875 186083 574941 186084
rect 574691 179212 574757 179213
rect 574691 179148 574692 179212
rect 574756 179148 574757 179212
rect 574691 179147 574757 179148
rect 567834 172938 567866 173494
rect 568422 172938 568454 173494
rect 567834 137494 568454 172938
rect 574691 171732 574757 171733
rect 574691 171668 574692 171732
rect 574756 171668 574757 171732
rect 574691 171667 574757 171668
rect 574694 152693 574754 171667
rect 574878 165885 574938 186083
rect 577794 183454 578414 218898
rect 577794 182898 577826 183454
rect 578382 182898 578414 183454
rect 574875 165884 574941 165885
rect 574875 165820 574876 165884
rect 574940 165820 574941 165884
rect 574875 165819 574941 165820
rect 574875 157316 574941 157317
rect 574875 157252 574876 157316
rect 574940 157252 574941 157316
rect 574875 157251 574941 157252
rect 574691 152692 574757 152693
rect 574691 152628 574692 152692
rect 574756 152628 574757 152692
rect 574691 152627 574757 152628
rect 569168 147454 569488 147486
rect 569168 147218 569210 147454
rect 569446 147218 569488 147454
rect 569168 147134 569488 147218
rect 569168 146898 569210 147134
rect 569446 146898 569488 147134
rect 569168 146866 569488 146898
rect 574691 142900 574757 142901
rect 574691 142836 574692 142900
rect 574756 142836 574757 142900
rect 574691 142835 574757 142836
rect 567834 136938 567866 137494
rect 568422 136938 568454 137494
rect 567834 101494 568454 136938
rect 574694 126037 574754 142835
rect 574878 139365 574938 157251
rect 577794 147454 578414 182898
rect 577794 146898 577826 147454
rect 578382 146898 578414 147454
rect 574875 139364 574941 139365
rect 574875 139300 574876 139364
rect 574940 139300 574941 139364
rect 574875 139299 574941 139300
rect 574875 128484 574941 128485
rect 574875 128420 574876 128484
rect 574940 128420 574941 128484
rect 574875 128419 574941 128420
rect 574691 126036 574757 126037
rect 574691 125972 574692 126036
rect 574756 125972 574757 126036
rect 574691 125971 574757 125972
rect 574691 114068 574757 114069
rect 574691 114004 574692 114068
rect 574756 114004 574757 114068
rect 574691 114003 574757 114004
rect 569168 111454 569488 111486
rect 569168 111218 569210 111454
rect 569446 111218 569488 111454
rect 569168 111134 569488 111218
rect 569168 110898 569210 111134
rect 569446 110898 569488 111134
rect 569168 110866 569488 110898
rect 567834 100938 567866 101494
rect 568422 100938 568454 101494
rect 567834 65494 568454 100938
rect 574694 99517 574754 114003
rect 574878 112845 574938 128419
rect 574875 112844 574941 112845
rect 574875 112780 574876 112844
rect 574940 112780 574941 112844
rect 574875 112779 574941 112780
rect 577794 111454 578414 146898
rect 577794 110898 577826 111454
rect 578382 110898 578414 111454
rect 574875 99652 574941 99653
rect 574875 99588 574876 99652
rect 574940 99588 574941 99652
rect 574875 99587 574941 99588
rect 574691 99516 574757 99517
rect 574691 99452 574692 99516
rect 574756 99452 574757 99516
rect 574691 99451 574757 99452
rect 574878 86189 574938 99587
rect 574875 86188 574941 86189
rect 574875 86124 574876 86188
rect 574940 86124 574941 86188
rect 574875 86123 574941 86124
rect 574691 85236 574757 85237
rect 574691 85172 574692 85236
rect 574756 85172 574757 85236
rect 574691 85171 574757 85172
rect 569168 75454 569488 75486
rect 569168 75218 569210 75454
rect 569446 75218 569488 75454
rect 569168 75134 569488 75218
rect 569168 74898 569210 75134
rect 569446 74898 569488 75134
rect 569168 74866 569488 74898
rect 574694 72997 574754 85171
rect 577794 75454 578414 110898
rect 577794 74898 577826 75454
rect 578382 74898 578414 75454
rect 574691 72996 574757 72997
rect 574691 72932 574692 72996
rect 574756 72932 574757 72996
rect 574691 72931 574757 72932
rect 574691 70820 574757 70821
rect 574691 70756 574692 70820
rect 574756 70756 574757 70820
rect 574691 70755 574757 70756
rect 567834 64938 567866 65494
rect 568422 64938 568454 65494
rect 567834 29494 568454 64938
rect 574694 59669 574754 70755
rect 574691 59668 574757 59669
rect 574691 59604 574692 59668
rect 574756 59604 574757 59668
rect 574691 59603 574757 59604
rect 574691 56404 574757 56405
rect 574691 56340 574692 56404
rect 574756 56340 574757 56404
rect 574691 56339 574757 56340
rect 574694 46341 574754 56339
rect 574691 46340 574757 46341
rect 574691 46276 574692 46340
rect 574756 46276 574757 46340
rect 574691 46275 574757 46276
rect 574691 41988 574757 41989
rect 574691 41924 574692 41988
rect 574756 41924 574757 41988
rect 574691 41923 574757 41924
rect 569168 39454 569488 39486
rect 569168 39218 569210 39454
rect 569446 39218 569488 39454
rect 569168 39134 569488 39218
rect 569168 38898 569210 39134
rect 569446 38898 569488 39134
rect 569168 38866 569488 38898
rect 574694 33149 574754 41923
rect 577794 39454 578414 74898
rect 577794 38898 577826 39454
rect 578382 38898 578414 39454
rect 574691 33148 574757 33149
rect 574691 33084 574692 33148
rect 574756 33084 574757 33148
rect 574691 33083 574757 33084
rect 567834 28938 567866 29494
rect 568422 28938 568454 29494
rect 567834 -7066 568454 28938
rect 575427 27572 575493 27573
rect 575427 27508 575428 27572
rect 575492 27508 575493 27572
rect 575427 27507 575493 27508
rect 575430 19821 575490 27507
rect 575427 19820 575493 19821
rect 575427 19756 575428 19820
rect 575492 19756 575493 19820
rect 575427 19755 575493 19756
rect 574691 13156 574757 13157
rect 574691 13092 574692 13156
rect 574756 13092 574757 13156
rect 574691 13091 574757 13092
rect 574694 6629 574754 13091
rect 574691 6628 574757 6629
rect 574691 6564 574692 6628
rect 574756 6564 574757 6628
rect 574691 6563 574757 6564
rect 567834 -7622 567866 -7066
rect 568422 -7622 568454 -7066
rect 567834 -7654 568454 -7622
rect 577794 3454 578414 38898
rect 577794 2898 577826 3454
rect 578382 2898 578414 3454
rect 577794 -346 578414 2898
rect 577794 -902 577826 -346
rect 578382 -902 578414 -346
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711002 592062 711558
rect 592618 711002 592650 711558
rect 591070 710598 591690 710630
rect 591070 710042 591102 710598
rect 591658 710042 591690 710598
rect 590110 709638 590730 709670
rect 590110 709082 590142 709638
rect 590698 709082 590730 709638
rect 589150 708678 589770 708710
rect 589150 708122 589182 708678
rect 589738 708122 589770 708678
rect 588190 707718 588810 707750
rect 588190 707162 588222 707718
rect 588778 707162 588810 707718
rect 587230 706758 587850 706790
rect 587230 706202 587262 706758
rect 587818 706202 587850 706758
rect 581514 705242 581546 705798
rect 582102 705242 582134 705798
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705242 586302 705798
rect 586858 705242 586890 705798
rect 581514 690618 581546 691174
rect 582102 690618 582134 691174
rect 581514 655174 582134 690618
rect 581514 654618 581546 655174
rect 582102 654618 582134 655174
rect 581514 619174 582134 654618
rect 581514 618618 581546 619174
rect 582102 618618 582134 619174
rect 581514 583174 582134 618618
rect 581514 582618 581546 583174
rect 582102 582618 582134 583174
rect 581514 547174 582134 582618
rect 581514 546618 581546 547174
rect 582102 546618 582134 547174
rect 581514 511174 582134 546618
rect 581514 510618 581546 511174
rect 582102 510618 582134 511174
rect 581514 475174 582134 510618
rect 581514 474618 581546 475174
rect 582102 474618 582134 475174
rect 581514 439174 582134 474618
rect 581514 438618 581546 439174
rect 582102 438618 582134 439174
rect 581514 403174 582134 438618
rect 581514 402618 581546 403174
rect 582102 402618 582134 403174
rect 581514 367174 582134 402618
rect 581514 366618 581546 367174
rect 582102 366618 582134 367174
rect 581514 331174 582134 366618
rect 581514 330618 581546 331174
rect 582102 330618 582134 331174
rect 581514 295174 582134 330618
rect 581514 294618 581546 295174
rect 582102 294618 582134 295174
rect 581514 259174 582134 294618
rect 581514 258618 581546 259174
rect 582102 258618 582134 259174
rect 581514 223174 582134 258618
rect 581514 222618 581546 223174
rect 582102 222618 582134 223174
rect 581514 187174 582134 222618
rect 581514 186618 581546 187174
rect 582102 186618 582134 187174
rect 581514 151174 582134 186618
rect 581514 150618 581546 151174
rect 582102 150618 582134 151174
rect 581514 115174 582134 150618
rect 581514 114618 581546 115174
rect 582102 114618 582134 115174
rect 581514 79174 582134 114618
rect 581514 78618 581546 79174
rect 582102 78618 582134 79174
rect 581514 43174 582134 78618
rect 581514 42618 581546 43174
rect 582102 42618 582134 43174
rect 581514 7174 582134 42618
rect 581514 6618 581546 7174
rect 582102 6618 582134 7174
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704282 585342 704838
rect 585898 704282 585930 704838
rect 585310 687454 585930 704282
rect 585310 686898 585342 687454
rect 585898 686898 585930 687454
rect 585310 651454 585930 686898
rect 585310 650898 585342 651454
rect 585898 650898 585930 651454
rect 585310 615454 585930 650898
rect 585310 614898 585342 615454
rect 585898 614898 585930 615454
rect 585310 579454 585930 614898
rect 585310 578898 585342 579454
rect 585898 578898 585930 579454
rect 585310 543454 585930 578898
rect 585310 542898 585342 543454
rect 585898 542898 585930 543454
rect 585310 507454 585930 542898
rect 585310 506898 585342 507454
rect 585898 506898 585930 507454
rect 585310 471454 585930 506898
rect 585310 470898 585342 471454
rect 585898 470898 585930 471454
rect 585310 435454 585930 470898
rect 585310 434898 585342 435454
rect 585898 434898 585930 435454
rect 585310 399454 585930 434898
rect 585310 398898 585342 399454
rect 585898 398898 585930 399454
rect 585310 363454 585930 398898
rect 585310 362898 585342 363454
rect 585898 362898 585930 363454
rect 585310 327454 585930 362898
rect 585310 326898 585342 327454
rect 585898 326898 585930 327454
rect 585310 291454 585930 326898
rect 585310 290898 585342 291454
rect 585898 290898 585930 291454
rect 585310 255454 585930 290898
rect 585310 254898 585342 255454
rect 585898 254898 585930 255454
rect 585310 219454 585930 254898
rect 585310 218898 585342 219454
rect 585898 218898 585930 219454
rect 585310 183454 585930 218898
rect 585310 182898 585342 183454
rect 585898 182898 585930 183454
rect 585310 147454 585930 182898
rect 585310 146898 585342 147454
rect 585898 146898 585930 147454
rect 585310 111454 585930 146898
rect 585310 110898 585342 111454
rect 585898 110898 585930 111454
rect 585310 75454 585930 110898
rect 585310 74898 585342 75454
rect 585898 74898 585930 75454
rect 585310 39454 585930 74898
rect 585310 38898 585342 39454
rect 585898 38898 585930 39454
rect 585310 3454 585930 38898
rect 585310 2898 585342 3454
rect 585898 2898 585930 3454
rect 585310 -346 585930 2898
rect 585310 -902 585342 -346
rect 585898 -902 585930 -346
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690618 586302 691174
rect 586858 690618 586890 691174
rect 586270 655174 586890 690618
rect 586270 654618 586302 655174
rect 586858 654618 586890 655174
rect 586270 619174 586890 654618
rect 586270 618618 586302 619174
rect 586858 618618 586890 619174
rect 586270 583174 586890 618618
rect 586270 582618 586302 583174
rect 586858 582618 586890 583174
rect 586270 547174 586890 582618
rect 586270 546618 586302 547174
rect 586858 546618 586890 547174
rect 586270 511174 586890 546618
rect 586270 510618 586302 511174
rect 586858 510618 586890 511174
rect 586270 475174 586890 510618
rect 586270 474618 586302 475174
rect 586858 474618 586890 475174
rect 586270 439174 586890 474618
rect 586270 438618 586302 439174
rect 586858 438618 586890 439174
rect 586270 403174 586890 438618
rect 586270 402618 586302 403174
rect 586858 402618 586890 403174
rect 586270 367174 586890 402618
rect 586270 366618 586302 367174
rect 586858 366618 586890 367174
rect 586270 331174 586890 366618
rect 586270 330618 586302 331174
rect 586858 330618 586890 331174
rect 586270 295174 586890 330618
rect 586270 294618 586302 295174
rect 586858 294618 586890 295174
rect 586270 259174 586890 294618
rect 586270 258618 586302 259174
rect 586858 258618 586890 259174
rect 586270 223174 586890 258618
rect 586270 222618 586302 223174
rect 586858 222618 586890 223174
rect 586270 187174 586890 222618
rect 586270 186618 586302 187174
rect 586858 186618 586890 187174
rect 586270 151174 586890 186618
rect 586270 150618 586302 151174
rect 586858 150618 586890 151174
rect 586270 115174 586890 150618
rect 586270 114618 586302 115174
rect 586858 114618 586890 115174
rect 586270 79174 586890 114618
rect 586270 78618 586302 79174
rect 586858 78618 586890 79174
rect 586270 43174 586890 78618
rect 586270 42618 586302 43174
rect 586858 42618 586890 43174
rect 586270 7174 586890 42618
rect 586270 6618 586302 7174
rect 586858 6618 586890 7174
rect 581514 -1862 581546 -1306
rect 582102 -1862 582134 -1306
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694338 587262 694894
rect 587818 694338 587850 694894
rect 587230 658894 587850 694338
rect 587230 658338 587262 658894
rect 587818 658338 587850 658894
rect 587230 622894 587850 658338
rect 587230 622338 587262 622894
rect 587818 622338 587850 622894
rect 587230 586894 587850 622338
rect 587230 586338 587262 586894
rect 587818 586338 587850 586894
rect 587230 550894 587850 586338
rect 587230 550338 587262 550894
rect 587818 550338 587850 550894
rect 587230 514894 587850 550338
rect 587230 514338 587262 514894
rect 587818 514338 587850 514894
rect 587230 478894 587850 514338
rect 587230 478338 587262 478894
rect 587818 478338 587850 478894
rect 587230 442894 587850 478338
rect 587230 442338 587262 442894
rect 587818 442338 587850 442894
rect 587230 406894 587850 442338
rect 587230 406338 587262 406894
rect 587818 406338 587850 406894
rect 587230 370894 587850 406338
rect 587230 370338 587262 370894
rect 587818 370338 587850 370894
rect 587230 334894 587850 370338
rect 587230 334338 587262 334894
rect 587818 334338 587850 334894
rect 587230 298894 587850 334338
rect 587230 298338 587262 298894
rect 587818 298338 587850 298894
rect 587230 262894 587850 298338
rect 587230 262338 587262 262894
rect 587818 262338 587850 262894
rect 587230 226894 587850 262338
rect 587230 226338 587262 226894
rect 587818 226338 587850 226894
rect 587230 190894 587850 226338
rect 587230 190338 587262 190894
rect 587818 190338 587850 190894
rect 587230 154894 587850 190338
rect 587230 154338 587262 154894
rect 587818 154338 587850 154894
rect 587230 118894 587850 154338
rect 587230 118338 587262 118894
rect 587818 118338 587850 118894
rect 587230 82894 587850 118338
rect 587230 82338 587262 82894
rect 587818 82338 587850 82894
rect 587230 46894 587850 82338
rect 587230 46338 587262 46894
rect 587818 46338 587850 46894
rect 587230 10894 587850 46338
rect 587230 10338 587262 10894
rect 587818 10338 587850 10894
rect 587230 -2266 587850 10338
rect 587230 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698058 588222 698614
rect 588778 698058 588810 698614
rect 588190 662614 588810 698058
rect 588190 662058 588222 662614
rect 588778 662058 588810 662614
rect 588190 626614 588810 662058
rect 588190 626058 588222 626614
rect 588778 626058 588810 626614
rect 588190 590614 588810 626058
rect 588190 590058 588222 590614
rect 588778 590058 588810 590614
rect 588190 554614 588810 590058
rect 588190 554058 588222 554614
rect 588778 554058 588810 554614
rect 588190 518614 588810 554058
rect 588190 518058 588222 518614
rect 588778 518058 588810 518614
rect 588190 482614 588810 518058
rect 588190 482058 588222 482614
rect 588778 482058 588810 482614
rect 588190 446614 588810 482058
rect 588190 446058 588222 446614
rect 588778 446058 588810 446614
rect 588190 410614 588810 446058
rect 588190 410058 588222 410614
rect 588778 410058 588810 410614
rect 588190 374614 588810 410058
rect 588190 374058 588222 374614
rect 588778 374058 588810 374614
rect 588190 338614 588810 374058
rect 588190 338058 588222 338614
rect 588778 338058 588810 338614
rect 588190 302614 588810 338058
rect 588190 302058 588222 302614
rect 588778 302058 588810 302614
rect 588190 266614 588810 302058
rect 588190 266058 588222 266614
rect 588778 266058 588810 266614
rect 588190 230614 588810 266058
rect 588190 230058 588222 230614
rect 588778 230058 588810 230614
rect 588190 194614 588810 230058
rect 588190 194058 588222 194614
rect 588778 194058 588810 194614
rect 588190 158614 588810 194058
rect 588190 158058 588222 158614
rect 588778 158058 588810 158614
rect 588190 122614 588810 158058
rect 588190 122058 588222 122614
rect 588778 122058 588810 122614
rect 588190 86614 588810 122058
rect 588190 86058 588222 86614
rect 588778 86058 588810 86614
rect 588190 50614 588810 86058
rect 588190 50058 588222 50614
rect 588778 50058 588810 50614
rect 588190 14614 588810 50058
rect 588190 14058 588222 14614
rect 588778 14058 588810 14614
rect 588190 -3226 588810 14058
rect 588190 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 665778 589182 666334
rect 589738 665778 589770 666334
rect 589150 630334 589770 665778
rect 589150 629778 589182 630334
rect 589738 629778 589770 630334
rect 589150 594334 589770 629778
rect 589150 593778 589182 594334
rect 589738 593778 589770 594334
rect 589150 558334 589770 593778
rect 589150 557778 589182 558334
rect 589738 557778 589770 558334
rect 589150 522334 589770 557778
rect 589150 521778 589182 522334
rect 589738 521778 589770 522334
rect 589150 486334 589770 521778
rect 589150 485778 589182 486334
rect 589738 485778 589770 486334
rect 589150 450334 589770 485778
rect 589150 449778 589182 450334
rect 589738 449778 589770 450334
rect 589150 414334 589770 449778
rect 589150 413778 589182 414334
rect 589738 413778 589770 414334
rect 589150 378334 589770 413778
rect 589150 377778 589182 378334
rect 589738 377778 589770 378334
rect 589150 342334 589770 377778
rect 589150 341778 589182 342334
rect 589738 341778 589770 342334
rect 589150 306334 589770 341778
rect 589150 305778 589182 306334
rect 589738 305778 589770 306334
rect 589150 270334 589770 305778
rect 589150 269778 589182 270334
rect 589738 269778 589770 270334
rect 589150 234334 589770 269778
rect 589150 233778 589182 234334
rect 589738 233778 589770 234334
rect 589150 198334 589770 233778
rect 589150 197778 589182 198334
rect 589738 197778 589770 198334
rect 589150 162334 589770 197778
rect 589150 161778 589182 162334
rect 589738 161778 589770 162334
rect 589150 126334 589770 161778
rect 589150 125778 589182 126334
rect 589738 125778 589770 126334
rect 589150 90334 589770 125778
rect 589150 89778 589182 90334
rect 589738 89778 589770 90334
rect 589150 54334 589770 89778
rect 589150 53778 589182 54334
rect 589738 53778 589770 54334
rect 589150 18334 589770 53778
rect 589150 17778 589182 18334
rect 589738 17778 589770 18334
rect 589150 -4186 589770 17778
rect 589150 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669498 590142 670054
rect 590698 669498 590730 670054
rect 590110 634054 590730 669498
rect 590110 633498 590142 634054
rect 590698 633498 590730 634054
rect 590110 598054 590730 633498
rect 590110 597498 590142 598054
rect 590698 597498 590730 598054
rect 590110 562054 590730 597498
rect 590110 561498 590142 562054
rect 590698 561498 590730 562054
rect 590110 526054 590730 561498
rect 590110 525498 590142 526054
rect 590698 525498 590730 526054
rect 590110 490054 590730 525498
rect 590110 489498 590142 490054
rect 590698 489498 590730 490054
rect 590110 454054 590730 489498
rect 590110 453498 590142 454054
rect 590698 453498 590730 454054
rect 590110 418054 590730 453498
rect 590110 417498 590142 418054
rect 590698 417498 590730 418054
rect 590110 382054 590730 417498
rect 590110 381498 590142 382054
rect 590698 381498 590730 382054
rect 590110 346054 590730 381498
rect 590110 345498 590142 346054
rect 590698 345498 590730 346054
rect 590110 310054 590730 345498
rect 590110 309498 590142 310054
rect 590698 309498 590730 310054
rect 590110 274054 590730 309498
rect 590110 273498 590142 274054
rect 590698 273498 590730 274054
rect 590110 238054 590730 273498
rect 590110 237498 590142 238054
rect 590698 237498 590730 238054
rect 590110 202054 590730 237498
rect 590110 201498 590142 202054
rect 590698 201498 590730 202054
rect 590110 166054 590730 201498
rect 590110 165498 590142 166054
rect 590698 165498 590730 166054
rect 590110 130054 590730 165498
rect 590110 129498 590142 130054
rect 590698 129498 590730 130054
rect 590110 94054 590730 129498
rect 590110 93498 590142 94054
rect 590698 93498 590730 94054
rect 590110 58054 590730 93498
rect 590110 57498 590142 58054
rect 590698 57498 590730 58054
rect 590110 22054 590730 57498
rect 590110 21498 590142 22054
rect 590698 21498 590730 22054
rect 590110 -5146 590730 21498
rect 590110 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673218 591102 673774
rect 591658 673218 591690 673774
rect 591070 637774 591690 673218
rect 591070 637218 591102 637774
rect 591658 637218 591690 637774
rect 591070 601774 591690 637218
rect 591070 601218 591102 601774
rect 591658 601218 591690 601774
rect 591070 565774 591690 601218
rect 591070 565218 591102 565774
rect 591658 565218 591690 565774
rect 591070 529774 591690 565218
rect 591070 529218 591102 529774
rect 591658 529218 591690 529774
rect 591070 493774 591690 529218
rect 591070 493218 591102 493774
rect 591658 493218 591690 493774
rect 591070 457774 591690 493218
rect 591070 457218 591102 457774
rect 591658 457218 591690 457774
rect 591070 421774 591690 457218
rect 591070 421218 591102 421774
rect 591658 421218 591690 421774
rect 591070 385774 591690 421218
rect 591070 385218 591102 385774
rect 591658 385218 591690 385774
rect 591070 349774 591690 385218
rect 591070 349218 591102 349774
rect 591658 349218 591690 349774
rect 591070 313774 591690 349218
rect 591070 313218 591102 313774
rect 591658 313218 591690 313774
rect 591070 277774 591690 313218
rect 591070 277218 591102 277774
rect 591658 277218 591690 277774
rect 591070 241774 591690 277218
rect 591070 241218 591102 241774
rect 591658 241218 591690 241774
rect 591070 205774 591690 241218
rect 591070 205218 591102 205774
rect 591658 205218 591690 205774
rect 591070 169774 591690 205218
rect 591070 169218 591102 169774
rect 591658 169218 591690 169774
rect 591070 133774 591690 169218
rect 591070 133218 591102 133774
rect 591658 133218 591690 133774
rect 591070 97774 591690 133218
rect 591070 97218 591102 97774
rect 591658 97218 591690 97774
rect 591070 61774 591690 97218
rect 591070 61218 591102 61774
rect 591658 61218 591690 61774
rect 591070 25774 591690 61218
rect 591070 25218 591102 25774
rect 591658 25218 591690 25774
rect 591070 -6106 591690 25218
rect 591070 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 676938 592062 677494
rect 592618 676938 592650 677494
rect 592030 641494 592650 676938
rect 592030 640938 592062 641494
rect 592618 640938 592650 641494
rect 592030 605494 592650 640938
rect 592030 604938 592062 605494
rect 592618 604938 592650 605494
rect 592030 569494 592650 604938
rect 592030 568938 592062 569494
rect 592618 568938 592650 569494
rect 592030 533494 592650 568938
rect 592030 532938 592062 533494
rect 592618 532938 592650 533494
rect 592030 497494 592650 532938
rect 592030 496938 592062 497494
rect 592618 496938 592650 497494
rect 592030 461494 592650 496938
rect 592030 460938 592062 461494
rect 592618 460938 592650 461494
rect 592030 425494 592650 460938
rect 592030 424938 592062 425494
rect 592618 424938 592650 425494
rect 592030 389494 592650 424938
rect 592030 388938 592062 389494
rect 592618 388938 592650 389494
rect 592030 353494 592650 388938
rect 592030 352938 592062 353494
rect 592618 352938 592650 353494
rect 592030 317494 592650 352938
rect 592030 316938 592062 317494
rect 592618 316938 592650 317494
rect 592030 281494 592650 316938
rect 592030 280938 592062 281494
rect 592618 280938 592650 281494
rect 592030 245494 592650 280938
rect 592030 244938 592062 245494
rect 592618 244938 592650 245494
rect 592030 209494 592650 244938
rect 592030 208938 592062 209494
rect 592618 208938 592650 209494
rect 592030 173494 592650 208938
rect 592030 172938 592062 173494
rect 592618 172938 592650 173494
rect 592030 137494 592650 172938
rect 592030 136938 592062 137494
rect 592618 136938 592650 137494
rect 592030 101494 592650 136938
rect 592030 100938 592062 101494
rect 592618 100938 592650 101494
rect 592030 65494 592650 100938
rect 592030 64938 592062 65494
rect 592618 64938 592650 65494
rect 592030 29494 592650 64938
rect 592030 28938 592062 29494
rect 592618 28938 592650 29494
rect 592030 -7066 592650 28938
rect 592030 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711002 -8138 711558
rect -8694 676938 -8138 677494
rect -8694 640938 -8138 641494
rect -8694 604938 -8138 605494
rect -8694 568938 -8138 569494
rect -8694 532938 -8138 533494
rect -8694 496938 -8138 497494
rect -8694 460938 -8138 461494
rect -8694 424938 -8138 425494
rect -8694 388938 -8138 389494
rect -8694 352938 -8138 353494
rect -8694 316938 -8138 317494
rect -8694 280938 -8138 281494
rect -8694 244938 -8138 245494
rect -8694 208938 -8138 209494
rect -8694 172938 -8138 173494
rect -8694 136938 -8138 137494
rect -8694 100938 -8138 101494
rect -8694 64938 -8138 65494
rect -8694 28938 -8138 29494
rect -7734 710042 -7178 710598
rect -7734 673218 -7178 673774
rect -7734 637218 -7178 637774
rect -7734 601218 -7178 601774
rect -7734 565218 -7178 565774
rect -7734 529218 -7178 529774
rect -7734 493218 -7178 493774
rect -7734 457218 -7178 457774
rect -7734 421218 -7178 421774
rect -7734 385218 -7178 385774
rect -7734 349218 -7178 349774
rect -7734 313218 -7178 313774
rect -7734 277218 -7178 277774
rect -7734 241218 -7178 241774
rect -7734 205218 -7178 205774
rect -7734 169218 -7178 169774
rect -7734 133218 -7178 133774
rect -7734 97218 -7178 97774
rect -7734 61218 -7178 61774
rect -7734 25218 -7178 25774
rect -6774 709082 -6218 709638
rect -6774 669498 -6218 670054
rect -6774 633498 -6218 634054
rect -6774 597498 -6218 598054
rect -6774 561498 -6218 562054
rect -6774 525498 -6218 526054
rect -6774 489498 -6218 490054
rect -6774 453498 -6218 454054
rect -6774 417498 -6218 418054
rect -6774 381498 -6218 382054
rect -6774 345498 -6218 346054
rect -6774 309498 -6218 310054
rect -6774 273498 -6218 274054
rect -6774 237498 -6218 238054
rect -6774 201498 -6218 202054
rect -6774 165498 -6218 166054
rect -6774 129498 -6218 130054
rect -6774 93498 -6218 94054
rect -6774 57498 -6218 58054
rect -6774 21498 -6218 22054
rect -5814 708122 -5258 708678
rect -5814 665778 -5258 666334
rect -5814 629778 -5258 630334
rect -5814 593778 -5258 594334
rect -5814 557778 -5258 558334
rect -5814 521778 -5258 522334
rect -5814 485778 -5258 486334
rect -5814 449778 -5258 450334
rect -5814 413778 -5258 414334
rect -5814 377778 -5258 378334
rect -5814 341778 -5258 342334
rect -5814 305778 -5258 306334
rect -5814 269778 -5258 270334
rect -5814 233778 -5258 234334
rect -5814 197778 -5258 198334
rect -5814 161778 -5258 162334
rect -5814 125778 -5258 126334
rect -5814 89778 -5258 90334
rect -5814 53778 -5258 54334
rect -5814 17778 -5258 18334
rect -4854 707162 -4298 707718
rect -4854 698058 -4298 698614
rect -4854 662058 -4298 662614
rect -4854 626058 -4298 626614
rect -4854 590058 -4298 590614
rect -4854 554058 -4298 554614
rect -4854 518058 -4298 518614
rect -4854 482058 -4298 482614
rect -4854 446058 -4298 446614
rect -4854 410058 -4298 410614
rect -4854 374058 -4298 374614
rect -4854 338058 -4298 338614
rect -4854 302058 -4298 302614
rect -4854 266058 -4298 266614
rect -4854 230058 -4298 230614
rect -4854 194058 -4298 194614
rect -4854 158058 -4298 158614
rect -4854 122058 -4298 122614
rect -4854 86058 -4298 86614
rect -4854 50058 -4298 50614
rect -4854 14058 -4298 14614
rect -3894 706202 -3338 706758
rect -3894 694338 -3338 694894
rect -3894 658338 -3338 658894
rect -3894 622338 -3338 622894
rect -3894 586338 -3338 586894
rect -3894 550338 -3338 550894
rect -3894 514338 -3338 514894
rect -3894 478338 -3338 478894
rect -3894 442338 -3338 442894
rect -3894 406338 -3338 406894
rect -3894 370338 -3338 370894
rect -3894 334338 -3338 334894
rect -3894 298338 -3338 298894
rect -3894 262338 -3338 262894
rect -3894 226338 -3338 226894
rect -3894 190338 -3338 190894
rect -3894 154338 -3338 154894
rect -3894 118338 -3338 118894
rect -3894 82338 -3338 82894
rect -3894 46338 -3338 46894
rect -3894 10338 -3338 10894
rect -2934 705242 -2378 705798
rect -2934 690618 -2378 691174
rect -2934 654618 -2378 655174
rect -2934 618618 -2378 619174
rect -2934 582618 -2378 583174
rect -2934 546618 -2378 547174
rect -2934 510618 -2378 511174
rect -2934 474618 -2378 475174
rect -2934 438618 -2378 439174
rect -2934 402618 -2378 403174
rect -2934 366618 -2378 367174
rect -2934 330618 -2378 331174
rect -2934 294618 -2378 295174
rect -2934 258618 -2378 259174
rect -2934 222618 -2378 223174
rect -2934 186618 -2378 187174
rect -2934 150618 -2378 151174
rect -2934 114618 -2378 115174
rect -2934 78618 -2378 79174
rect -2934 42618 -2378 43174
rect -2934 6618 -2378 7174
rect -1974 704282 -1418 704838
rect -1974 686898 -1418 687454
rect -1974 650898 -1418 651454
rect -1974 614898 -1418 615454
rect -1974 578898 -1418 579454
rect -1974 542898 -1418 543454
rect -1974 506898 -1418 507454
rect -1974 470898 -1418 471454
rect -1974 434898 -1418 435454
rect -1974 398898 -1418 399454
rect -1974 362898 -1418 363454
rect -1974 326898 -1418 327454
rect -1974 290898 -1418 291454
rect -1974 254898 -1418 255454
rect -1974 218898 -1418 219454
rect -1974 182898 -1418 183454
rect -1974 146898 -1418 147454
rect -1974 110898 -1418 111454
rect -1974 74898 -1418 75454
rect -1974 38898 -1418 39454
rect -1974 2898 -1418 3454
rect -1974 -902 -1418 -346
rect 1826 704282 2382 704838
rect 1826 686898 2382 687454
rect 1826 650898 2382 651454
rect 1826 614898 2382 615454
rect 1826 578898 2382 579454
rect 1826 542898 2382 543454
rect 1826 506898 2382 507454
rect 1826 470898 2382 471454
rect 1826 434898 2382 435454
rect 1826 398898 2382 399454
rect 5546 705242 6102 705798
rect 5546 690618 6102 691174
rect 5546 654618 6102 655174
rect 5546 618618 6102 619174
rect 5546 582618 6102 583174
rect 5546 546618 6102 547174
rect 5546 510618 6102 511174
rect 5546 474618 6102 475174
rect 5546 438618 6102 439174
rect 5546 402618 6102 403174
rect 1826 362898 2382 363454
rect 1826 326898 2382 327454
rect 5546 366618 6102 367174
rect 5546 330618 6102 331174
rect 1826 290898 2382 291454
rect 5546 294618 6102 295174
rect 1826 254898 2382 255454
rect 1826 218898 2382 219454
rect 1826 182898 2382 183454
rect 1826 146898 2382 147454
rect 9266 706202 9822 706758
rect 9266 694338 9822 694894
rect 9266 658338 9822 658894
rect 9266 622338 9822 622894
rect 9266 586338 9822 586894
rect 9266 550338 9822 550894
rect 9266 514338 9822 514894
rect 9266 478338 9822 478894
rect 9266 442338 9822 442894
rect 9266 406338 9822 406894
rect 9266 370338 9822 370894
rect 9266 334338 9822 334894
rect 9266 298338 9822 298894
rect 5546 258618 6102 259174
rect 9266 262338 9822 262894
rect 5546 222618 6102 223174
rect 9266 226338 9822 226894
rect 9266 190338 9822 190894
rect 5546 186618 6102 187174
rect 5546 150618 6102 151174
rect 1826 110898 2382 111454
rect 9266 154338 9822 154894
rect 5546 114618 6102 115174
rect 1826 74898 2382 75454
rect 1826 38898 2382 39454
rect 1826 2898 2382 3454
rect 1826 -902 2382 -346
rect -2934 -1862 -2378 -1306
rect -3894 -2822 -3338 -2266
rect -4854 -3782 -4298 -3226
rect -5814 -4742 -5258 -4186
rect -6774 -5702 -6218 -5146
rect -7734 -6662 -7178 -6106
rect -8694 -7622 -8138 -7066
rect 9266 118338 9822 118894
rect 5546 78618 6102 79174
rect 9266 82338 9822 82894
rect 9266 46338 9822 46894
rect 5546 42618 6102 43174
rect 5546 6618 6102 7174
rect 9266 10338 9822 10894
rect 5546 -1862 6102 -1306
rect 9266 -2822 9822 -2266
rect 12986 707162 13542 707718
rect 12986 698058 13542 698614
rect 12986 662058 13542 662614
rect 12986 626058 13542 626614
rect 12986 590058 13542 590614
rect 12986 554058 13542 554614
rect 12986 518058 13542 518614
rect 12986 482058 13542 482614
rect 12986 446058 13542 446614
rect 12986 410058 13542 410614
rect 12986 374058 13542 374614
rect 12986 338058 13542 338614
rect 16706 708122 17262 708678
rect 16706 665778 17262 666334
rect 16706 629778 17262 630334
rect 16706 593778 17262 594334
rect 16706 557778 17262 558334
rect 16706 521778 17262 522334
rect 16706 485778 17262 486334
rect 16706 449778 17262 450334
rect 16706 413778 17262 414334
rect 16706 377778 17262 378334
rect 16706 341778 17262 342334
rect 16250 327218 16486 327454
rect 16250 326898 16486 327134
rect 12986 302058 13542 302614
rect 16706 305778 17262 306334
rect 16250 291218 16486 291454
rect 16250 290898 16486 291134
rect 12986 266058 13542 266614
rect 16706 269778 17262 270334
rect 16250 255218 16486 255454
rect 16250 254898 16486 255134
rect 12986 230058 13542 230614
rect 16706 233778 17262 234334
rect 16250 219218 16486 219454
rect 16250 218898 16486 219134
rect 12986 194058 13542 194614
rect 16706 197778 17262 198334
rect 16250 183218 16486 183454
rect 16250 182898 16486 183134
rect 12986 158058 13542 158614
rect 16706 161778 17262 162334
rect 16250 147218 16486 147454
rect 16250 146898 16486 147134
rect 12986 122058 13542 122614
rect 16706 125778 17262 126334
rect 16250 111218 16486 111454
rect 16250 110898 16486 111134
rect 12986 86058 13542 86614
rect 16706 89778 17262 90334
rect 16250 75218 16486 75454
rect 16250 74898 16486 75134
rect 12986 50058 13542 50614
rect 16706 53778 17262 54334
rect 16250 39218 16486 39454
rect 16250 38898 16486 39134
rect 12986 14058 13542 14614
rect 12986 -3782 13542 -3226
rect 16706 17778 17262 18334
rect 16706 -4742 17262 -4186
rect 20426 709082 20982 709638
rect 20426 669498 20982 670054
rect 20426 633498 20982 634054
rect 20426 597498 20982 598054
rect 20426 561498 20982 562054
rect 20426 525498 20982 526054
rect 20426 489498 20982 490054
rect 20426 453498 20982 454054
rect 20426 417498 20982 418054
rect 20426 381498 20982 382054
rect 20426 345498 20982 346054
rect 20426 309498 20982 310054
rect 20426 273498 20982 274054
rect 20426 237498 20982 238054
rect 20426 201498 20982 202054
rect 20426 165498 20982 166054
rect 20426 129498 20982 130054
rect 20426 93498 20982 94054
rect 20426 57498 20982 58054
rect 20426 21498 20982 22054
rect 20426 -5702 20982 -5146
rect 24146 710042 24702 710598
rect 24146 673218 24702 673774
rect 24146 637218 24702 637774
rect 24146 601218 24702 601774
rect 24146 565218 24702 565774
rect 24146 529218 24702 529774
rect 24146 493218 24702 493774
rect 24146 457218 24702 457774
rect 24146 421218 24702 421774
rect 24146 385218 24702 385774
rect 24146 349218 24702 349774
rect 24146 313218 24702 313774
rect 24146 277218 24702 277774
rect 24146 241218 24702 241774
rect 24146 205218 24702 205774
rect 24146 169218 24702 169774
rect 24146 133218 24702 133774
rect 24146 97218 24702 97774
rect 24146 61218 24702 61774
rect 24146 25218 24702 25774
rect 24146 -6662 24702 -6106
rect 27866 711002 28422 711558
rect 27866 676938 28422 677494
rect 27866 640938 28422 641494
rect 27866 604938 28422 605494
rect 27866 568938 28422 569494
rect 27866 532938 28422 533494
rect 27866 496938 28422 497494
rect 27866 460938 28422 461494
rect 27866 424938 28422 425494
rect 27866 388938 28422 389494
rect 27866 352938 28422 353494
rect 37826 704282 38382 704838
rect 37826 686898 38382 687454
rect 37826 650898 38382 651454
rect 37826 614898 38382 615454
rect 37826 578898 38382 579454
rect 37826 542898 38382 543454
rect 37826 506898 38382 507454
rect 37826 470898 38382 471454
rect 37826 434898 38382 435454
rect 37826 398898 38382 399454
rect 37826 362898 38382 363454
rect 31610 330938 31846 331174
rect 31610 330618 31846 330854
rect 27866 316938 28422 317494
rect 37826 326898 38382 327454
rect 31610 294938 31846 295174
rect 31610 294618 31846 294854
rect 27866 280938 28422 281494
rect 37826 290898 38382 291454
rect 31610 258938 31846 259174
rect 31610 258618 31846 258854
rect 27866 244938 28422 245494
rect 37826 254898 38382 255454
rect 31610 222938 31846 223174
rect 31610 222618 31846 222854
rect 27866 208938 28422 209494
rect 37826 218898 38382 219454
rect 31610 186938 31846 187174
rect 31610 186618 31846 186854
rect 27866 172938 28422 173494
rect 37826 182898 38382 183454
rect 31610 150938 31846 151174
rect 31610 150618 31846 150854
rect 27866 136938 28422 137494
rect 37826 146898 38382 147454
rect 31610 114938 31846 115174
rect 31610 114618 31846 114854
rect 27866 100938 28422 101494
rect 37826 110898 38382 111454
rect 31610 78938 31846 79174
rect 31610 78618 31846 78854
rect 27866 64938 28422 65494
rect 37826 74898 38382 75454
rect 31610 42938 31846 43174
rect 31610 42618 31846 42854
rect 27866 28938 28422 29494
rect 37826 38898 38382 39454
rect 31610 6938 31846 7174
rect 31610 6618 31846 6854
rect 37826 2898 38382 3454
rect 27866 -7622 28422 -7066
rect 37826 -902 38382 -346
rect 41546 705242 42102 705798
rect 41546 690618 42102 691174
rect 41546 654618 42102 655174
rect 41546 618618 42102 619174
rect 41546 582618 42102 583174
rect 41546 546618 42102 547174
rect 41546 510618 42102 511174
rect 41546 474618 42102 475174
rect 41546 438618 42102 439174
rect 41546 402618 42102 403174
rect 41546 366618 42102 367174
rect 41546 330618 42102 331174
rect 41546 294618 42102 295174
rect 41546 258618 42102 259174
rect 41546 222618 42102 223174
rect 41546 186618 42102 187174
rect 41546 150618 42102 151174
rect 41546 114618 42102 115174
rect 41546 78618 42102 79174
rect 41546 42618 42102 43174
rect 41546 6618 42102 7174
rect 41546 -1862 42102 -1306
rect 45266 706202 45822 706758
rect 45266 694338 45822 694894
rect 45266 658338 45822 658894
rect 45266 622338 45822 622894
rect 45266 586338 45822 586894
rect 45266 550338 45822 550894
rect 45266 514338 45822 514894
rect 45266 478338 45822 478894
rect 45266 442338 45822 442894
rect 45266 406338 45822 406894
rect 45266 370338 45822 370894
rect 45266 334338 45822 334894
rect 48986 707162 49542 707718
rect 48986 698058 49542 698614
rect 48986 662058 49542 662614
rect 48986 626058 49542 626614
rect 48986 590058 49542 590614
rect 48986 554058 49542 554614
rect 48986 518058 49542 518614
rect 48986 482058 49542 482614
rect 48986 446058 49542 446614
rect 48986 410058 49542 410614
rect 48986 374058 49542 374614
rect 48986 338058 49542 338614
rect 46970 327218 47206 327454
rect 46970 326898 47206 327134
rect 45266 298338 45822 298894
rect 48986 302058 49542 302614
rect 46970 291218 47206 291454
rect 46970 290898 47206 291134
rect 45266 262338 45822 262894
rect 48986 266058 49542 266614
rect 46970 255218 47206 255454
rect 46970 254898 47206 255134
rect 45266 226338 45822 226894
rect 48986 230058 49542 230614
rect 46970 219218 47206 219454
rect 46970 218898 47206 219134
rect 45266 190338 45822 190894
rect 48986 194058 49542 194614
rect 46970 183218 47206 183454
rect 46970 182898 47206 183134
rect 45266 154338 45822 154894
rect 48986 158058 49542 158614
rect 46970 147218 47206 147454
rect 46970 146898 47206 147134
rect 45266 118338 45822 118894
rect 48986 122058 49542 122614
rect 46970 111218 47206 111454
rect 46970 110898 47206 111134
rect 45266 82338 45822 82894
rect 48986 86058 49542 86614
rect 46970 75218 47206 75454
rect 46970 74898 47206 75134
rect 45266 46338 45822 46894
rect 48986 50058 49542 50614
rect 46970 39218 47206 39454
rect 46970 38898 47206 39134
rect 45266 10338 45822 10894
rect 48986 14058 49542 14614
rect 45266 -2822 45822 -2266
rect 48986 -3782 49542 -3226
rect 52706 708122 53262 708678
rect 52706 665778 53262 666334
rect 52706 629778 53262 630334
rect 52706 593778 53262 594334
rect 52706 557778 53262 558334
rect 52706 521778 53262 522334
rect 52706 485778 53262 486334
rect 52706 449778 53262 450334
rect 52706 413778 53262 414334
rect 52706 377778 53262 378334
rect 52706 341778 53262 342334
rect 52706 305778 53262 306334
rect 52706 269778 53262 270334
rect 52706 233778 53262 234334
rect 52706 197778 53262 198334
rect 52706 161778 53262 162334
rect 52706 125778 53262 126334
rect 52706 89778 53262 90334
rect 52706 53778 53262 54334
rect 52706 17778 53262 18334
rect 52706 -4742 53262 -4186
rect 56426 709082 56982 709638
rect 56426 669498 56982 670054
rect 56426 633498 56982 634054
rect 56426 597498 56982 598054
rect 56426 561498 56982 562054
rect 56426 525498 56982 526054
rect 56426 489498 56982 490054
rect 56426 453498 56982 454054
rect 56426 417498 56982 418054
rect 56426 381498 56982 382054
rect 56426 345498 56982 346054
rect 56426 309498 56982 310054
rect 56426 273498 56982 274054
rect 56426 237498 56982 238054
rect 56426 201498 56982 202054
rect 56426 165498 56982 166054
rect 56426 129498 56982 130054
rect 56426 93498 56982 94054
rect 56426 57498 56982 58054
rect 56426 21498 56982 22054
rect 60146 710042 60702 710598
rect 60146 673218 60702 673774
rect 60146 637218 60702 637774
rect 60146 601218 60702 601774
rect 60146 565218 60702 565774
rect 60146 529218 60702 529774
rect 60146 493218 60702 493774
rect 60146 457218 60702 457774
rect 60146 421218 60702 421774
rect 60146 385218 60702 385774
rect 60146 349218 60702 349774
rect 63866 711002 64422 711558
rect 63866 676938 64422 677494
rect 63866 640938 64422 641494
rect 63866 604938 64422 605494
rect 63866 568938 64422 569494
rect 63866 532938 64422 533494
rect 63866 496938 64422 497494
rect 63866 460938 64422 461494
rect 63866 424938 64422 425494
rect 63866 388938 64422 389494
rect 63866 352938 64422 353494
rect 62330 330938 62566 331174
rect 62330 330618 62566 330854
rect 60146 313218 60702 313774
rect 63866 316938 64422 317494
rect 62330 294938 62566 295174
rect 62330 294618 62566 294854
rect 60146 277218 60702 277774
rect 63866 280938 64422 281494
rect 62330 258938 62566 259174
rect 62330 258618 62566 258854
rect 60146 241218 60702 241774
rect 63866 244938 64422 245494
rect 62330 222938 62566 223174
rect 62330 222618 62566 222854
rect 60146 205218 60702 205774
rect 63866 208938 64422 209494
rect 62330 186938 62566 187174
rect 62330 186618 62566 186854
rect 60146 169218 60702 169774
rect 63866 172938 64422 173494
rect 62330 150938 62566 151174
rect 62330 150618 62566 150854
rect 60146 133218 60702 133774
rect 63866 136938 64422 137494
rect 62330 114938 62566 115174
rect 62330 114618 62566 114854
rect 60146 97218 60702 97774
rect 63866 100938 64422 101494
rect 62330 78938 62566 79174
rect 62330 78618 62566 78854
rect 60146 61218 60702 61774
rect 63866 64938 64422 65494
rect 62330 42938 62566 43174
rect 62330 42618 62566 42854
rect 60146 25218 60702 25774
rect 56426 -5702 56982 -5146
rect 63866 28938 64422 29494
rect 62330 6938 62566 7174
rect 62330 6618 62566 6854
rect 60146 -6662 60702 -6106
rect 63866 -7622 64422 -7066
rect 73826 704282 74382 704838
rect 73826 686898 74382 687454
rect 73826 650898 74382 651454
rect 73826 614898 74382 615454
rect 73826 578898 74382 579454
rect 73826 542898 74382 543454
rect 73826 506898 74382 507454
rect 73826 470898 74382 471454
rect 73826 434898 74382 435454
rect 73826 398898 74382 399454
rect 73826 362898 74382 363454
rect 77546 705242 78102 705798
rect 77546 690618 78102 691174
rect 77546 654618 78102 655174
rect 77546 618618 78102 619174
rect 77546 582618 78102 583174
rect 77546 546618 78102 547174
rect 77546 510618 78102 511174
rect 77546 474618 78102 475174
rect 77546 438618 78102 439174
rect 77546 402618 78102 403174
rect 77546 366618 78102 367174
rect 81266 706202 81822 706758
rect 81266 694338 81822 694894
rect 81266 658338 81822 658894
rect 81266 622338 81822 622894
rect 81266 586338 81822 586894
rect 81266 550338 81822 550894
rect 81266 514338 81822 514894
rect 81266 478338 81822 478894
rect 81266 442338 81822 442894
rect 81266 406338 81822 406894
rect 81266 370338 81822 370894
rect 81266 334338 81822 334894
rect 73826 326898 74382 327454
rect 77690 327218 77926 327454
rect 77690 326898 77926 327134
rect 81266 298338 81822 298894
rect 73826 290898 74382 291454
rect 77690 291218 77926 291454
rect 77690 290898 77926 291134
rect 81266 262338 81822 262894
rect 73826 254898 74382 255454
rect 77690 255218 77926 255454
rect 77690 254898 77926 255134
rect 81266 226338 81822 226894
rect 73826 218898 74382 219454
rect 77690 219218 77926 219454
rect 77690 218898 77926 219134
rect 81266 190338 81822 190894
rect 73826 182898 74382 183454
rect 77690 183218 77926 183454
rect 77690 182898 77926 183134
rect 81266 154338 81822 154894
rect 73826 146898 74382 147454
rect 77690 147218 77926 147454
rect 77690 146898 77926 147134
rect 81266 118338 81822 118894
rect 73826 110898 74382 111454
rect 77690 111218 77926 111454
rect 77690 110898 77926 111134
rect 81266 82338 81822 82894
rect 73826 74898 74382 75454
rect 77690 75218 77926 75454
rect 77690 74898 77926 75134
rect 81266 46338 81822 46894
rect 73826 38898 74382 39454
rect 77690 39218 77926 39454
rect 77690 38898 77926 39134
rect 73826 2898 74382 3454
rect 73826 -902 74382 -346
rect 81266 10338 81822 10894
rect 81266 -2822 81822 -2266
rect 84986 707162 85542 707718
rect 84986 698058 85542 698614
rect 84986 662058 85542 662614
rect 84986 626058 85542 626614
rect 84986 590058 85542 590614
rect 84986 554058 85542 554614
rect 84986 518058 85542 518614
rect 84986 482058 85542 482614
rect 84986 446058 85542 446614
rect 84986 410058 85542 410614
rect 84986 374058 85542 374614
rect 84986 338058 85542 338614
rect 84986 302058 85542 302614
rect 84986 266058 85542 266614
rect 84986 230058 85542 230614
rect 84986 194058 85542 194614
rect 84986 158058 85542 158614
rect 84986 122058 85542 122614
rect 84986 86058 85542 86614
rect 84986 50058 85542 50614
rect 84986 14058 85542 14614
rect 84986 -3782 85542 -3226
rect 88706 708122 89262 708678
rect 88706 665778 89262 666334
rect 88706 629778 89262 630334
rect 88706 593778 89262 594334
rect 88706 557778 89262 558334
rect 88706 521778 89262 522334
rect 88706 485778 89262 486334
rect 88706 449778 89262 450334
rect 88706 413778 89262 414334
rect 88706 377778 89262 378334
rect 92426 709082 92982 709638
rect 92426 669498 92982 670054
rect 92426 633498 92982 634054
rect 92426 597498 92982 598054
rect 92426 561498 92982 562054
rect 92426 525498 92982 526054
rect 92426 489498 92982 490054
rect 92426 453498 92982 454054
rect 92426 417498 92982 418054
rect 92426 381498 92982 382054
rect 96146 710042 96702 710598
rect 96146 673218 96702 673774
rect 96146 637218 96702 637774
rect 96146 601218 96702 601774
rect 96146 565218 96702 565774
rect 96146 529218 96702 529774
rect 96146 493218 96702 493774
rect 96146 457218 96702 457774
rect 96146 421218 96702 421774
rect 96146 385218 96702 385774
rect 88706 341778 89262 342334
rect 96146 349218 96702 349774
rect 93050 330938 93286 331174
rect 93050 330618 93286 330854
rect 88706 305778 89262 306334
rect 96146 313218 96702 313774
rect 93050 294938 93286 295174
rect 93050 294618 93286 294854
rect 88706 269778 89262 270334
rect 96146 277218 96702 277774
rect 93050 258938 93286 259174
rect 93050 258618 93286 258854
rect 88706 233778 89262 234334
rect 96146 241218 96702 241774
rect 93050 222938 93286 223174
rect 93050 222618 93286 222854
rect 88706 197778 89262 198334
rect 96146 205218 96702 205774
rect 93050 186938 93286 187174
rect 93050 186618 93286 186854
rect 88706 161778 89262 162334
rect 96146 169218 96702 169774
rect 93050 150938 93286 151174
rect 93050 150618 93286 150854
rect 88706 125778 89262 126334
rect 96146 133218 96702 133774
rect 93050 114938 93286 115174
rect 93050 114618 93286 114854
rect 88706 89778 89262 90334
rect 96146 97218 96702 97774
rect 93050 78938 93286 79174
rect 93050 78618 93286 78854
rect 88706 53778 89262 54334
rect 96146 61218 96702 61774
rect 93050 42938 93286 43174
rect 93050 42618 93286 42854
rect 88706 17778 89262 18334
rect 96146 25218 96702 25774
rect 93050 6938 93286 7174
rect 93050 6618 93286 6854
rect 88706 -4742 89262 -4186
rect 96146 -6662 96702 -6106
rect 99866 711002 100422 711558
rect 99866 676938 100422 677494
rect 99866 640938 100422 641494
rect 99866 604938 100422 605494
rect 99866 568938 100422 569494
rect 99866 532938 100422 533494
rect 99866 496938 100422 497494
rect 99866 460938 100422 461494
rect 99866 424938 100422 425494
rect 99866 388938 100422 389494
rect 99866 352938 100422 353494
rect 109826 704282 110382 704838
rect 109826 686898 110382 687454
rect 109826 650898 110382 651454
rect 109826 614898 110382 615454
rect 109826 578898 110382 579454
rect 109826 542898 110382 543454
rect 109826 506898 110382 507454
rect 109826 470898 110382 471454
rect 109826 434898 110382 435454
rect 109826 398898 110382 399454
rect 109826 362898 110382 363454
rect 108410 327218 108646 327454
rect 108410 326898 108646 327134
rect 109826 326898 110382 327454
rect 99866 316938 100422 317494
rect 108410 291218 108646 291454
rect 108410 290898 108646 291134
rect 109826 290898 110382 291454
rect 99866 280938 100422 281494
rect 108410 255218 108646 255454
rect 108410 254898 108646 255134
rect 109826 254898 110382 255454
rect 99866 244938 100422 245494
rect 108410 219218 108646 219454
rect 108410 218898 108646 219134
rect 109826 218898 110382 219454
rect 99866 208938 100422 209494
rect 108410 183218 108646 183454
rect 108410 182898 108646 183134
rect 109826 182898 110382 183454
rect 99866 172938 100422 173494
rect 108410 147218 108646 147454
rect 108410 146898 108646 147134
rect 109826 146898 110382 147454
rect 99866 136938 100422 137494
rect 108410 111218 108646 111454
rect 108410 110898 108646 111134
rect 109826 110898 110382 111454
rect 99866 100938 100422 101494
rect 108410 75218 108646 75454
rect 108410 74898 108646 75134
rect 109826 74898 110382 75454
rect 99866 64938 100422 65494
rect 108410 39218 108646 39454
rect 108410 38898 108646 39134
rect 109826 38898 110382 39454
rect 99866 28938 100422 29494
rect 99866 -7622 100422 -7066
rect 109826 2898 110382 3454
rect 109826 -902 110382 -346
rect 113546 705242 114102 705798
rect 113546 690618 114102 691174
rect 113546 654618 114102 655174
rect 113546 618618 114102 619174
rect 113546 582618 114102 583174
rect 113546 546618 114102 547174
rect 113546 510618 114102 511174
rect 113546 474618 114102 475174
rect 113546 438618 114102 439174
rect 113546 402618 114102 403174
rect 113546 366618 114102 367174
rect 113546 330618 114102 331174
rect 113546 294618 114102 295174
rect 113546 258618 114102 259174
rect 113546 222618 114102 223174
rect 113546 186618 114102 187174
rect 113546 150618 114102 151174
rect 113546 114618 114102 115174
rect 113546 78618 114102 79174
rect 113546 42618 114102 43174
rect 113546 6618 114102 7174
rect 113546 -1862 114102 -1306
rect 117266 706202 117822 706758
rect 117266 694338 117822 694894
rect 117266 658338 117822 658894
rect 117266 622338 117822 622894
rect 117266 586338 117822 586894
rect 117266 550338 117822 550894
rect 117266 514338 117822 514894
rect 117266 478338 117822 478894
rect 117266 442338 117822 442894
rect 117266 406338 117822 406894
rect 117266 370338 117822 370894
rect 117266 334338 117822 334894
rect 117266 298338 117822 298894
rect 117266 262338 117822 262894
rect 117266 226338 117822 226894
rect 117266 190338 117822 190894
rect 117266 154338 117822 154894
rect 117266 118338 117822 118894
rect 117266 82338 117822 82894
rect 117266 46338 117822 46894
rect 117266 10338 117822 10894
rect 117266 -2822 117822 -2266
rect 120986 707162 121542 707718
rect 120986 698058 121542 698614
rect 120986 662058 121542 662614
rect 120986 626058 121542 626614
rect 120986 590058 121542 590614
rect 120986 554058 121542 554614
rect 120986 518058 121542 518614
rect 120986 482058 121542 482614
rect 120986 446058 121542 446614
rect 120986 410058 121542 410614
rect 120986 374058 121542 374614
rect 120986 338058 121542 338614
rect 124706 708122 125262 708678
rect 124706 665778 125262 666334
rect 124706 629778 125262 630334
rect 124706 593778 125262 594334
rect 124706 557778 125262 558334
rect 124706 521778 125262 522334
rect 124706 485778 125262 486334
rect 124706 449778 125262 450334
rect 124706 413778 125262 414334
rect 124706 377778 125262 378334
rect 124706 341778 125262 342334
rect 123770 330938 124006 331174
rect 123770 330618 124006 330854
rect 120986 302058 121542 302614
rect 124706 305778 125262 306334
rect 123770 294938 124006 295174
rect 123770 294618 124006 294854
rect 120986 266058 121542 266614
rect 124706 269778 125262 270334
rect 123770 258938 124006 259174
rect 123770 258618 124006 258854
rect 120986 230058 121542 230614
rect 124706 233778 125262 234334
rect 123770 222938 124006 223174
rect 123770 222618 124006 222854
rect 120986 194058 121542 194614
rect 124706 197778 125262 198334
rect 123770 186938 124006 187174
rect 123770 186618 124006 186854
rect 120986 158058 121542 158614
rect 124706 161778 125262 162334
rect 123770 150938 124006 151174
rect 123770 150618 124006 150854
rect 120986 122058 121542 122614
rect 124706 125778 125262 126334
rect 123770 114938 124006 115174
rect 123770 114618 124006 114854
rect 120986 86058 121542 86614
rect 124706 89778 125262 90334
rect 123770 78938 124006 79174
rect 123770 78618 124006 78854
rect 120986 50058 121542 50614
rect 124706 53778 125262 54334
rect 123770 42938 124006 43174
rect 123770 42618 124006 42854
rect 120986 14058 121542 14614
rect 124706 17778 125262 18334
rect 123770 6938 124006 7174
rect 123770 6618 124006 6854
rect 120986 -3782 121542 -3226
rect 124706 -4742 125262 -4186
rect 128426 709082 128982 709638
rect 128426 669498 128982 670054
rect 128426 633498 128982 634054
rect 128426 597498 128982 598054
rect 128426 561498 128982 562054
rect 128426 525498 128982 526054
rect 128426 489498 128982 490054
rect 128426 453498 128982 454054
rect 128426 417498 128982 418054
rect 128426 381498 128982 382054
rect 128426 345498 128982 346054
rect 128426 309498 128982 310054
rect 128426 273498 128982 274054
rect 128426 237498 128982 238054
rect 128426 201498 128982 202054
rect 128426 165498 128982 166054
rect 128426 129498 128982 130054
rect 128426 93498 128982 94054
rect 128426 57498 128982 58054
rect 128426 21498 128982 22054
rect 128426 -5702 128982 -5146
rect 132146 710042 132702 710598
rect 132146 673218 132702 673774
rect 132146 637218 132702 637774
rect 132146 601218 132702 601774
rect 132146 565218 132702 565774
rect 132146 529218 132702 529774
rect 132146 493218 132702 493774
rect 132146 457218 132702 457774
rect 132146 421218 132702 421774
rect 132146 385218 132702 385774
rect 132146 349218 132702 349774
rect 132146 313218 132702 313774
rect 132146 277218 132702 277774
rect 132146 241218 132702 241774
rect 132146 205218 132702 205774
rect 132146 169218 132702 169774
rect 132146 133218 132702 133774
rect 132146 97218 132702 97774
rect 132146 61218 132702 61774
rect 132146 25218 132702 25774
rect 132146 -6662 132702 -6106
rect 135866 711002 136422 711558
rect 135866 676938 136422 677494
rect 135866 640938 136422 641494
rect 135866 604938 136422 605494
rect 135866 568938 136422 569494
rect 135866 532938 136422 533494
rect 135866 496938 136422 497494
rect 135866 460938 136422 461494
rect 135866 424938 136422 425494
rect 135866 388938 136422 389494
rect 135866 352938 136422 353494
rect 145826 704282 146382 704838
rect 145826 686898 146382 687454
rect 145826 650898 146382 651454
rect 145826 614898 146382 615454
rect 145826 578898 146382 579454
rect 145826 542898 146382 543454
rect 145826 506898 146382 507454
rect 145826 470898 146382 471454
rect 145826 434898 146382 435454
rect 145826 398898 146382 399454
rect 145826 362898 146382 363454
rect 139130 327218 139366 327454
rect 139130 326898 139366 327134
rect 145826 326898 146382 327454
rect 135866 316938 136422 317494
rect 139130 291218 139366 291454
rect 139130 290898 139366 291134
rect 145826 290898 146382 291454
rect 135866 280938 136422 281494
rect 139130 255218 139366 255454
rect 139130 254898 139366 255134
rect 145826 254898 146382 255454
rect 135866 244938 136422 245494
rect 139130 219218 139366 219454
rect 139130 218898 139366 219134
rect 145826 218898 146382 219454
rect 135866 208938 136422 209494
rect 139130 183218 139366 183454
rect 139130 182898 139366 183134
rect 145826 182898 146382 183454
rect 135866 172938 136422 173494
rect 139130 147218 139366 147454
rect 139130 146898 139366 147134
rect 145826 146898 146382 147454
rect 135866 136938 136422 137494
rect 139130 111218 139366 111454
rect 139130 110898 139366 111134
rect 145826 110898 146382 111454
rect 135866 100938 136422 101494
rect 139130 75218 139366 75454
rect 139130 74898 139366 75134
rect 145826 74898 146382 75454
rect 135866 64938 136422 65494
rect 139130 39218 139366 39454
rect 139130 38898 139366 39134
rect 145826 38898 146382 39454
rect 135866 28938 136422 29494
rect 135866 -7622 136422 -7066
rect 145826 2898 146382 3454
rect 145826 -902 146382 -346
rect 149546 705242 150102 705798
rect 149546 690618 150102 691174
rect 149546 654618 150102 655174
rect 149546 618618 150102 619174
rect 149546 582618 150102 583174
rect 149546 546618 150102 547174
rect 149546 510618 150102 511174
rect 149546 474618 150102 475174
rect 149546 438618 150102 439174
rect 149546 402618 150102 403174
rect 149546 366618 150102 367174
rect 149546 330618 150102 331174
rect 149546 294618 150102 295174
rect 149546 258618 150102 259174
rect 149546 222618 150102 223174
rect 149546 186618 150102 187174
rect 149546 150618 150102 151174
rect 149546 114618 150102 115174
rect 149546 78618 150102 79174
rect 149546 42618 150102 43174
rect 149546 6618 150102 7174
rect 149546 -1862 150102 -1306
rect 153266 706202 153822 706758
rect 153266 694338 153822 694894
rect 153266 658338 153822 658894
rect 153266 622338 153822 622894
rect 153266 586338 153822 586894
rect 153266 550338 153822 550894
rect 153266 514338 153822 514894
rect 153266 478338 153822 478894
rect 153266 442338 153822 442894
rect 153266 406338 153822 406894
rect 153266 370338 153822 370894
rect 153266 334338 153822 334894
rect 156986 707162 157542 707718
rect 156986 698058 157542 698614
rect 156986 662058 157542 662614
rect 156986 626058 157542 626614
rect 156986 590058 157542 590614
rect 156986 554058 157542 554614
rect 156986 518058 157542 518614
rect 156986 482058 157542 482614
rect 156986 446058 157542 446614
rect 156986 410058 157542 410614
rect 156986 374058 157542 374614
rect 156986 338058 157542 338614
rect 154490 330938 154726 331174
rect 154490 330618 154726 330854
rect 153266 298338 153822 298894
rect 156986 302058 157542 302614
rect 154490 294938 154726 295174
rect 154490 294618 154726 294854
rect 153266 262338 153822 262894
rect 156986 266058 157542 266614
rect 154490 258938 154726 259174
rect 154490 258618 154726 258854
rect 153266 226338 153822 226894
rect 156986 230058 157542 230614
rect 154490 222938 154726 223174
rect 154490 222618 154726 222854
rect 153266 190338 153822 190894
rect 156986 194058 157542 194614
rect 154490 186938 154726 187174
rect 154490 186618 154726 186854
rect 153266 154338 153822 154894
rect 156986 158058 157542 158614
rect 154490 150938 154726 151174
rect 154490 150618 154726 150854
rect 153266 118338 153822 118894
rect 156986 122058 157542 122614
rect 154490 114938 154726 115174
rect 154490 114618 154726 114854
rect 153266 82338 153822 82894
rect 156986 86058 157542 86614
rect 154490 78938 154726 79174
rect 154490 78618 154726 78854
rect 153266 46338 153822 46894
rect 156986 50058 157542 50614
rect 154490 42938 154726 43174
rect 154490 42618 154726 42854
rect 153266 10338 153822 10894
rect 156986 14058 157542 14614
rect 154490 6938 154726 7174
rect 154490 6618 154726 6854
rect 153266 -2822 153822 -2266
rect 156986 -3782 157542 -3226
rect 160706 708122 161262 708678
rect 160706 665778 161262 666334
rect 160706 629778 161262 630334
rect 160706 593778 161262 594334
rect 160706 557778 161262 558334
rect 160706 521778 161262 522334
rect 160706 485778 161262 486334
rect 160706 449778 161262 450334
rect 160706 413778 161262 414334
rect 160706 377778 161262 378334
rect 160706 341778 161262 342334
rect 160706 305778 161262 306334
rect 160706 269778 161262 270334
rect 160706 233778 161262 234334
rect 160706 197778 161262 198334
rect 160706 161778 161262 162334
rect 160706 125778 161262 126334
rect 160706 89778 161262 90334
rect 160706 53778 161262 54334
rect 160706 17778 161262 18334
rect 160706 -4742 161262 -4186
rect 164426 709082 164982 709638
rect 164426 669498 164982 670054
rect 164426 633498 164982 634054
rect 164426 597498 164982 598054
rect 164426 561498 164982 562054
rect 164426 525498 164982 526054
rect 164426 489498 164982 490054
rect 164426 453498 164982 454054
rect 164426 417498 164982 418054
rect 164426 381498 164982 382054
rect 164426 345498 164982 346054
rect 164426 309498 164982 310054
rect 164426 273498 164982 274054
rect 164426 237498 164982 238054
rect 164426 201498 164982 202054
rect 164426 165498 164982 166054
rect 164426 129498 164982 130054
rect 164426 93498 164982 94054
rect 164426 57498 164982 58054
rect 164426 21498 164982 22054
rect 164426 -5702 164982 -5146
rect 168146 710042 168702 710598
rect 168146 673218 168702 673774
rect 168146 637218 168702 637774
rect 168146 601218 168702 601774
rect 168146 565218 168702 565774
rect 168146 529218 168702 529774
rect 168146 493218 168702 493774
rect 168146 457218 168702 457774
rect 168146 421218 168702 421774
rect 168146 385218 168702 385774
rect 168146 349218 168702 349774
rect 171866 711002 172422 711558
rect 171866 676938 172422 677494
rect 171866 640938 172422 641494
rect 171866 604938 172422 605494
rect 171866 568938 172422 569494
rect 171866 532938 172422 533494
rect 171866 496938 172422 497494
rect 171866 460938 172422 461494
rect 171866 424938 172422 425494
rect 171866 388938 172422 389494
rect 171866 352938 172422 353494
rect 169850 327218 170086 327454
rect 169850 326898 170086 327134
rect 168146 313218 168702 313774
rect 171866 316938 172422 317494
rect 169850 291218 170086 291454
rect 169850 290898 170086 291134
rect 168146 277218 168702 277774
rect 171866 280938 172422 281494
rect 169850 255218 170086 255454
rect 169850 254898 170086 255134
rect 168146 241218 168702 241774
rect 171866 244938 172422 245494
rect 169850 219218 170086 219454
rect 169850 218898 170086 219134
rect 168146 205218 168702 205774
rect 171866 208938 172422 209494
rect 169850 183218 170086 183454
rect 169850 182898 170086 183134
rect 168146 169218 168702 169774
rect 171866 172938 172422 173494
rect 169850 147218 170086 147454
rect 169850 146898 170086 147134
rect 168146 133218 168702 133774
rect 171866 136938 172422 137494
rect 169850 111218 170086 111454
rect 169850 110898 170086 111134
rect 168146 97218 168702 97774
rect 171866 100938 172422 101494
rect 169850 75218 170086 75454
rect 169850 74898 170086 75134
rect 168146 61218 168702 61774
rect 171866 64938 172422 65494
rect 169850 39218 170086 39454
rect 169850 38898 170086 39134
rect 168146 25218 168702 25774
rect 168146 -6662 168702 -6106
rect 171866 28938 172422 29494
rect 171866 -7622 172422 -7066
rect 181826 704282 182382 704838
rect 181826 686898 182382 687454
rect 181826 650898 182382 651454
rect 181826 614898 182382 615454
rect 181826 578898 182382 579454
rect 181826 542898 182382 543454
rect 181826 506898 182382 507454
rect 181826 470898 182382 471454
rect 181826 434898 182382 435454
rect 181826 398898 182382 399454
rect 181826 362898 182382 363454
rect 185546 705242 186102 705798
rect 185546 690618 186102 691174
rect 185546 654618 186102 655174
rect 185546 618618 186102 619174
rect 185546 582618 186102 583174
rect 185546 546618 186102 547174
rect 185546 510618 186102 511174
rect 185546 474618 186102 475174
rect 185546 438618 186102 439174
rect 185546 402618 186102 403174
rect 185546 366618 186102 367174
rect 189266 706202 189822 706758
rect 189266 694338 189822 694894
rect 189266 658338 189822 658894
rect 189266 622338 189822 622894
rect 189266 586338 189822 586894
rect 189266 550338 189822 550894
rect 189266 514338 189822 514894
rect 189266 478338 189822 478894
rect 189266 442338 189822 442894
rect 189266 406338 189822 406894
rect 189266 370338 189822 370894
rect 189266 334338 189822 334894
rect 185210 330938 185446 331174
rect 185210 330618 185446 330854
rect 181826 326898 182382 327454
rect 189266 298338 189822 298894
rect 185210 294938 185446 295174
rect 185210 294618 185446 294854
rect 181826 290898 182382 291454
rect 189266 262338 189822 262894
rect 185210 258938 185446 259174
rect 185210 258618 185446 258854
rect 181826 254898 182382 255454
rect 189266 226338 189822 226894
rect 185210 222938 185446 223174
rect 185210 222618 185446 222854
rect 181826 218898 182382 219454
rect 189266 190338 189822 190894
rect 185210 186938 185446 187174
rect 185210 186618 185446 186854
rect 181826 182898 182382 183454
rect 189266 154338 189822 154894
rect 185210 150938 185446 151174
rect 185210 150618 185446 150854
rect 181826 146898 182382 147454
rect 189266 118338 189822 118894
rect 185210 114938 185446 115174
rect 185210 114618 185446 114854
rect 181826 110898 182382 111454
rect 189266 82338 189822 82894
rect 185210 78938 185446 79174
rect 185210 78618 185446 78854
rect 181826 74898 182382 75454
rect 189266 46338 189822 46894
rect 185210 42938 185446 43174
rect 185210 42618 185446 42854
rect 181826 38898 182382 39454
rect 189266 10338 189822 10894
rect 185210 6938 185446 7174
rect 185210 6618 185446 6854
rect 181826 2898 182382 3454
rect 181826 -902 182382 -346
rect 189266 -2822 189822 -2266
rect 192986 707162 193542 707718
rect 192986 698058 193542 698614
rect 192986 662058 193542 662614
rect 192986 626058 193542 626614
rect 192986 590058 193542 590614
rect 192986 554058 193542 554614
rect 192986 518058 193542 518614
rect 192986 482058 193542 482614
rect 192986 446058 193542 446614
rect 192986 410058 193542 410614
rect 192986 374058 193542 374614
rect 192986 338058 193542 338614
rect 192986 302058 193542 302614
rect 192986 266058 193542 266614
rect 192986 230058 193542 230614
rect 192986 194058 193542 194614
rect 192986 158058 193542 158614
rect 192986 122058 193542 122614
rect 192986 86058 193542 86614
rect 192986 50058 193542 50614
rect 192986 14058 193542 14614
rect 192986 -3782 193542 -3226
rect 196706 708122 197262 708678
rect 196706 665778 197262 666334
rect 196706 629778 197262 630334
rect 196706 593778 197262 594334
rect 196706 557778 197262 558334
rect 196706 521778 197262 522334
rect 196706 485778 197262 486334
rect 196706 449778 197262 450334
rect 196706 413778 197262 414334
rect 196706 377778 197262 378334
rect 200426 709082 200982 709638
rect 200426 669498 200982 670054
rect 200426 633498 200982 634054
rect 200426 597498 200982 598054
rect 200426 561498 200982 562054
rect 200426 525498 200982 526054
rect 200426 489498 200982 490054
rect 200426 453498 200982 454054
rect 200426 417498 200982 418054
rect 200426 381498 200982 382054
rect 204146 710042 204702 710598
rect 204146 673218 204702 673774
rect 204146 637218 204702 637774
rect 204146 601218 204702 601774
rect 204146 565218 204702 565774
rect 204146 529218 204702 529774
rect 204146 493218 204702 493774
rect 204146 457218 204702 457774
rect 204146 421218 204702 421774
rect 204146 385218 204702 385774
rect 196706 341778 197262 342334
rect 204146 349218 204702 349774
rect 200570 327218 200806 327454
rect 200570 326898 200806 327134
rect 196706 305778 197262 306334
rect 204146 313218 204702 313774
rect 200570 291218 200806 291454
rect 200570 290898 200806 291134
rect 196706 269778 197262 270334
rect 204146 277218 204702 277774
rect 200570 255218 200806 255454
rect 200570 254898 200806 255134
rect 196706 233778 197262 234334
rect 204146 241218 204702 241774
rect 200570 219218 200806 219454
rect 200570 218898 200806 219134
rect 196706 197778 197262 198334
rect 204146 205218 204702 205774
rect 200570 183218 200806 183454
rect 200570 182898 200806 183134
rect 196706 161778 197262 162334
rect 204146 169218 204702 169774
rect 200570 147218 200806 147454
rect 200570 146898 200806 147134
rect 196706 125778 197262 126334
rect 204146 133218 204702 133774
rect 200570 111218 200806 111454
rect 200570 110898 200806 111134
rect 196706 89778 197262 90334
rect 204146 97218 204702 97774
rect 200570 75218 200806 75454
rect 200570 74898 200806 75134
rect 196706 53778 197262 54334
rect 204146 61218 204702 61774
rect 200570 39218 200806 39454
rect 200570 38898 200806 39134
rect 196706 17778 197262 18334
rect 196706 -4742 197262 -4186
rect 204146 25218 204702 25774
rect 204146 -6662 204702 -6106
rect 207866 711002 208422 711558
rect 207866 676938 208422 677494
rect 207866 640938 208422 641494
rect 207866 604938 208422 605494
rect 207866 568938 208422 569494
rect 207866 532938 208422 533494
rect 207866 496938 208422 497494
rect 207866 460938 208422 461494
rect 207866 424938 208422 425494
rect 207866 388938 208422 389494
rect 207866 352938 208422 353494
rect 217826 704282 218382 704838
rect 217826 686898 218382 687454
rect 217826 650898 218382 651454
rect 217826 614898 218382 615454
rect 217826 578898 218382 579454
rect 217826 542898 218382 543454
rect 217826 506898 218382 507454
rect 217826 470898 218382 471454
rect 217826 434898 218382 435454
rect 217826 398898 218382 399454
rect 217826 362898 218382 363454
rect 215930 330938 216166 331174
rect 215930 330618 216166 330854
rect 207866 316938 208422 317494
rect 217826 326898 218382 327454
rect 215930 294938 216166 295174
rect 215930 294618 216166 294854
rect 207866 280938 208422 281494
rect 217826 290898 218382 291454
rect 215930 258938 216166 259174
rect 215930 258618 216166 258854
rect 207866 244938 208422 245494
rect 217826 254898 218382 255454
rect 215930 222938 216166 223174
rect 215930 222618 216166 222854
rect 207866 208938 208422 209494
rect 217826 218898 218382 219454
rect 215930 186938 216166 187174
rect 215930 186618 216166 186854
rect 207866 172938 208422 173494
rect 217826 182898 218382 183454
rect 215930 150938 216166 151174
rect 215930 150618 216166 150854
rect 207866 136938 208422 137494
rect 217826 146898 218382 147454
rect 215930 114938 216166 115174
rect 215930 114618 216166 114854
rect 207866 100938 208422 101494
rect 217826 110898 218382 111454
rect 215930 78938 216166 79174
rect 215930 78618 216166 78854
rect 207866 64938 208422 65494
rect 217826 74898 218382 75454
rect 215930 42938 216166 43174
rect 215930 42618 216166 42854
rect 207866 28938 208422 29494
rect 217826 38898 218382 39454
rect 215930 6938 216166 7174
rect 215930 6618 216166 6854
rect 207866 -7622 208422 -7066
rect 217826 2898 218382 3454
rect 217826 -902 218382 -346
rect 221546 705242 222102 705798
rect 221546 690618 222102 691174
rect 221546 654618 222102 655174
rect 221546 618618 222102 619174
rect 221546 582618 222102 583174
rect 221546 546618 222102 547174
rect 221546 510618 222102 511174
rect 221546 474618 222102 475174
rect 221546 438618 222102 439174
rect 221546 402618 222102 403174
rect 221546 366618 222102 367174
rect 221546 330618 222102 331174
rect 221546 294618 222102 295174
rect 221546 258618 222102 259174
rect 221546 222618 222102 223174
rect 221546 186618 222102 187174
rect 221546 150618 222102 151174
rect 221546 114618 222102 115174
rect 221546 78618 222102 79174
rect 221546 42618 222102 43174
rect 221546 6618 222102 7174
rect 221546 -1862 222102 -1306
rect 225266 706202 225822 706758
rect 225266 694338 225822 694894
rect 225266 658338 225822 658894
rect 225266 622338 225822 622894
rect 225266 586338 225822 586894
rect 225266 550338 225822 550894
rect 225266 514338 225822 514894
rect 225266 478338 225822 478894
rect 225266 442338 225822 442894
rect 225266 406338 225822 406894
rect 225266 370338 225822 370894
rect 225266 334338 225822 334894
rect 225266 298338 225822 298894
rect 225266 262338 225822 262894
rect 225266 226338 225822 226894
rect 225266 190338 225822 190894
rect 225266 154338 225822 154894
rect 225266 118338 225822 118894
rect 225266 82338 225822 82894
rect 225266 46338 225822 46894
rect 225266 10338 225822 10894
rect 225266 -2822 225822 -2266
rect 228986 707162 229542 707718
rect 228986 698058 229542 698614
rect 228986 662058 229542 662614
rect 228986 626058 229542 626614
rect 228986 590058 229542 590614
rect 228986 554058 229542 554614
rect 228986 518058 229542 518614
rect 228986 482058 229542 482614
rect 228986 446058 229542 446614
rect 228986 410058 229542 410614
rect 228986 374058 229542 374614
rect 228986 338058 229542 338614
rect 232706 708122 233262 708678
rect 232706 665778 233262 666334
rect 232706 629778 233262 630334
rect 232706 593778 233262 594334
rect 232706 557778 233262 558334
rect 232706 521778 233262 522334
rect 232706 485778 233262 486334
rect 232706 449778 233262 450334
rect 232706 413778 233262 414334
rect 232706 377778 233262 378334
rect 232706 341778 233262 342334
rect 231290 327218 231526 327454
rect 231290 326898 231526 327134
rect 228986 302058 229542 302614
rect 232706 305778 233262 306334
rect 231290 291218 231526 291454
rect 231290 290898 231526 291134
rect 228986 266058 229542 266614
rect 232706 269778 233262 270334
rect 231290 255218 231526 255454
rect 231290 254898 231526 255134
rect 228986 230058 229542 230614
rect 232706 233778 233262 234334
rect 231290 219218 231526 219454
rect 231290 218898 231526 219134
rect 228986 194058 229542 194614
rect 232706 197778 233262 198334
rect 231290 183218 231526 183454
rect 231290 182898 231526 183134
rect 228986 158058 229542 158614
rect 232706 161778 233262 162334
rect 231290 147218 231526 147454
rect 231290 146898 231526 147134
rect 228986 122058 229542 122614
rect 232706 125778 233262 126334
rect 231290 111218 231526 111454
rect 231290 110898 231526 111134
rect 228986 86058 229542 86614
rect 232706 89778 233262 90334
rect 231290 75218 231526 75454
rect 231290 74898 231526 75134
rect 228986 50058 229542 50614
rect 232706 53778 233262 54334
rect 231290 39218 231526 39454
rect 231290 38898 231526 39134
rect 228986 14058 229542 14614
rect 228986 -3782 229542 -3226
rect 232706 17778 233262 18334
rect 232706 -4742 233262 -4186
rect 236426 709082 236982 709638
rect 236426 669498 236982 670054
rect 236426 633498 236982 634054
rect 236426 597498 236982 598054
rect 236426 561498 236982 562054
rect 236426 525498 236982 526054
rect 236426 489498 236982 490054
rect 236426 453498 236982 454054
rect 236426 417498 236982 418054
rect 236426 381498 236982 382054
rect 236426 345498 236982 346054
rect 236426 309498 236982 310054
rect 236426 273498 236982 274054
rect 236426 237498 236982 238054
rect 236426 201498 236982 202054
rect 236426 165498 236982 166054
rect 236426 129498 236982 130054
rect 236426 93498 236982 94054
rect 236426 57498 236982 58054
rect 236426 21498 236982 22054
rect 236426 -5702 236982 -5146
rect 240146 710042 240702 710598
rect 240146 673218 240702 673774
rect 240146 637218 240702 637774
rect 240146 601218 240702 601774
rect 240146 565218 240702 565774
rect 240146 529218 240702 529774
rect 240146 493218 240702 493774
rect 240146 457218 240702 457774
rect 240146 421218 240702 421774
rect 240146 385218 240702 385774
rect 240146 349218 240702 349774
rect 240146 313218 240702 313774
rect 240146 277218 240702 277774
rect 240146 241218 240702 241774
rect 240146 205218 240702 205774
rect 240146 169218 240702 169774
rect 240146 133218 240702 133774
rect 240146 97218 240702 97774
rect 240146 61218 240702 61774
rect 240146 25218 240702 25774
rect 240146 -6662 240702 -6106
rect 243866 711002 244422 711558
rect 243866 676938 244422 677494
rect 243866 640938 244422 641494
rect 243866 604938 244422 605494
rect 243866 568938 244422 569494
rect 243866 532938 244422 533494
rect 243866 496938 244422 497494
rect 243866 460938 244422 461494
rect 243866 424938 244422 425494
rect 243866 388938 244422 389494
rect 243866 352938 244422 353494
rect 253826 704282 254382 704838
rect 253826 686898 254382 687454
rect 253826 650898 254382 651454
rect 253826 614898 254382 615454
rect 253826 578898 254382 579454
rect 253826 542898 254382 543454
rect 253826 506898 254382 507454
rect 253826 470898 254382 471454
rect 253826 434898 254382 435454
rect 253826 398898 254382 399454
rect 253826 362898 254382 363454
rect 246650 330938 246886 331174
rect 246650 330618 246886 330854
rect 243866 316938 244422 317494
rect 253826 326898 254382 327454
rect 246650 294938 246886 295174
rect 246650 294618 246886 294854
rect 243866 280938 244422 281494
rect 253826 290898 254382 291454
rect 246650 258938 246886 259174
rect 246650 258618 246886 258854
rect 243866 244938 244422 245494
rect 253826 254898 254382 255454
rect 246650 222938 246886 223174
rect 246650 222618 246886 222854
rect 243866 208938 244422 209494
rect 253826 218898 254382 219454
rect 246650 186938 246886 187174
rect 246650 186618 246886 186854
rect 243866 172938 244422 173494
rect 253826 182898 254382 183454
rect 246650 150938 246886 151174
rect 246650 150618 246886 150854
rect 243866 136938 244422 137494
rect 253826 146898 254382 147454
rect 246650 114938 246886 115174
rect 246650 114618 246886 114854
rect 243866 100938 244422 101494
rect 253826 110898 254382 111454
rect 246650 78938 246886 79174
rect 246650 78618 246886 78854
rect 243866 64938 244422 65494
rect 253826 74898 254382 75454
rect 246650 42938 246886 43174
rect 246650 42618 246886 42854
rect 243866 28938 244422 29494
rect 253826 38898 254382 39454
rect 246650 6938 246886 7174
rect 246650 6618 246886 6854
rect 243866 -7622 244422 -7066
rect 253826 2898 254382 3454
rect 253826 -902 254382 -346
rect 257546 705242 258102 705798
rect 257546 690618 258102 691174
rect 257546 654618 258102 655174
rect 257546 618618 258102 619174
rect 257546 582618 258102 583174
rect 257546 546618 258102 547174
rect 257546 510618 258102 511174
rect 257546 474618 258102 475174
rect 257546 438618 258102 439174
rect 257546 402618 258102 403174
rect 257546 366618 258102 367174
rect 261266 706202 261822 706758
rect 261266 694338 261822 694894
rect 261266 658338 261822 658894
rect 261266 622338 261822 622894
rect 261266 586338 261822 586894
rect 261266 550338 261822 550894
rect 261266 514338 261822 514894
rect 261266 478338 261822 478894
rect 261266 442338 261822 442894
rect 261266 406338 261822 406894
rect 261266 370338 261822 370894
rect 264986 707162 265542 707718
rect 264986 698058 265542 698614
rect 264986 662058 265542 662614
rect 264986 626058 265542 626614
rect 264986 590058 265542 590614
rect 264986 554058 265542 554614
rect 264986 518058 265542 518614
rect 264986 482058 265542 482614
rect 264986 446058 265542 446614
rect 264986 410058 265542 410614
rect 264986 374058 265542 374614
rect 257546 330618 258102 331174
rect 264986 338058 265542 338614
rect 262010 327218 262246 327454
rect 262010 326898 262246 327134
rect 257546 294618 258102 295174
rect 264986 302058 265542 302614
rect 262010 291218 262246 291454
rect 262010 290898 262246 291134
rect 257546 258618 258102 259174
rect 264986 266058 265542 266614
rect 262010 255218 262246 255454
rect 262010 254898 262246 255134
rect 257546 222618 258102 223174
rect 264986 230058 265542 230614
rect 262010 219218 262246 219454
rect 262010 218898 262246 219134
rect 257546 186618 258102 187174
rect 264986 194058 265542 194614
rect 262010 183218 262246 183454
rect 262010 182898 262246 183134
rect 257546 150618 258102 151174
rect 264986 158058 265542 158614
rect 262010 147218 262246 147454
rect 262010 146898 262246 147134
rect 257546 114618 258102 115174
rect 264986 122058 265542 122614
rect 262010 111218 262246 111454
rect 262010 110898 262246 111134
rect 257546 78618 258102 79174
rect 264986 86058 265542 86614
rect 262010 75218 262246 75454
rect 262010 74898 262246 75134
rect 257546 42618 258102 43174
rect 264986 50058 265542 50614
rect 262010 39218 262246 39454
rect 262010 38898 262246 39134
rect 257546 6618 258102 7174
rect 257546 -1862 258102 -1306
rect 264986 14058 265542 14614
rect 264986 -3782 265542 -3226
rect 268706 708122 269262 708678
rect 268706 665778 269262 666334
rect 268706 629778 269262 630334
rect 268706 593778 269262 594334
rect 268706 557778 269262 558334
rect 268706 521778 269262 522334
rect 268706 485778 269262 486334
rect 268706 449778 269262 450334
rect 268706 413778 269262 414334
rect 268706 377778 269262 378334
rect 268706 341778 269262 342334
rect 268706 305778 269262 306334
rect 268706 269778 269262 270334
rect 268706 233778 269262 234334
rect 268706 197778 269262 198334
rect 268706 161778 269262 162334
rect 268706 125778 269262 126334
rect 268706 89778 269262 90334
rect 268706 53778 269262 54334
rect 268706 17778 269262 18334
rect 268706 -4742 269262 -4186
rect 272426 709082 272982 709638
rect 272426 669498 272982 670054
rect 272426 633498 272982 634054
rect 272426 597498 272982 598054
rect 272426 561498 272982 562054
rect 272426 525498 272982 526054
rect 272426 489498 272982 490054
rect 272426 453498 272982 454054
rect 272426 417498 272982 418054
rect 272426 381498 272982 382054
rect 272426 345498 272982 346054
rect 272426 309498 272982 310054
rect 272426 273498 272982 274054
rect 272426 237498 272982 238054
rect 272426 201498 272982 202054
rect 272426 165498 272982 166054
rect 272426 129498 272982 130054
rect 272426 93498 272982 94054
rect 272426 57498 272982 58054
rect 272426 21498 272982 22054
rect 272426 -5702 272982 -5146
rect 276146 710042 276702 710598
rect 276146 673218 276702 673774
rect 276146 637218 276702 637774
rect 276146 601218 276702 601774
rect 276146 565218 276702 565774
rect 276146 529218 276702 529774
rect 276146 493218 276702 493774
rect 276146 457218 276702 457774
rect 276146 421218 276702 421774
rect 276146 385218 276702 385774
rect 276146 349218 276702 349774
rect 279866 711002 280422 711558
rect 279866 676938 280422 677494
rect 279866 640938 280422 641494
rect 279866 604938 280422 605494
rect 279866 568938 280422 569494
rect 279866 532938 280422 533494
rect 279866 496938 280422 497494
rect 279866 460938 280422 461494
rect 279866 424938 280422 425494
rect 279866 388938 280422 389494
rect 279866 352938 280422 353494
rect 277370 330938 277606 331174
rect 277370 330618 277606 330854
rect 276146 313218 276702 313774
rect 279866 316938 280422 317494
rect 277370 294938 277606 295174
rect 277370 294618 277606 294854
rect 276146 277218 276702 277774
rect 279866 280938 280422 281494
rect 277370 258938 277606 259174
rect 277370 258618 277606 258854
rect 276146 241218 276702 241774
rect 279866 244938 280422 245494
rect 277370 222938 277606 223174
rect 277370 222618 277606 222854
rect 276146 205218 276702 205774
rect 279866 208938 280422 209494
rect 277370 186938 277606 187174
rect 277370 186618 277606 186854
rect 276146 169218 276702 169774
rect 279866 172938 280422 173494
rect 277370 150938 277606 151174
rect 277370 150618 277606 150854
rect 276146 133218 276702 133774
rect 279866 136938 280422 137494
rect 277370 114938 277606 115174
rect 277370 114618 277606 114854
rect 276146 97218 276702 97774
rect 279866 100938 280422 101494
rect 277370 78938 277606 79174
rect 277370 78618 277606 78854
rect 276146 61218 276702 61774
rect 279866 64938 280422 65494
rect 277370 42938 277606 43174
rect 277370 42618 277606 42854
rect 276146 25218 276702 25774
rect 279866 28938 280422 29494
rect 277370 6938 277606 7174
rect 277370 6618 277606 6854
rect 276146 -6662 276702 -6106
rect 279866 -7622 280422 -7066
rect 289826 704282 290382 704838
rect 289826 686898 290382 687454
rect 289826 650898 290382 651454
rect 289826 614898 290382 615454
rect 289826 578898 290382 579454
rect 289826 542898 290382 543454
rect 289826 506898 290382 507454
rect 289826 470898 290382 471454
rect 289826 434898 290382 435454
rect 289826 398898 290382 399454
rect 289826 362898 290382 363454
rect 293546 705242 294102 705798
rect 293546 690618 294102 691174
rect 293546 654618 294102 655174
rect 293546 618618 294102 619174
rect 293546 582618 294102 583174
rect 293546 546618 294102 547174
rect 293546 510618 294102 511174
rect 293546 474618 294102 475174
rect 293546 438618 294102 439174
rect 293546 402618 294102 403174
rect 293546 366618 294102 367174
rect 293546 330618 294102 331174
rect 289826 326898 290382 327454
rect 292730 327218 292966 327454
rect 292730 326898 292966 327134
rect 293546 294618 294102 295174
rect 289826 290898 290382 291454
rect 292730 291218 292966 291454
rect 292730 290898 292966 291134
rect 293546 258618 294102 259174
rect 289826 254898 290382 255454
rect 292730 255218 292966 255454
rect 292730 254898 292966 255134
rect 293546 222618 294102 223174
rect 289826 218898 290382 219454
rect 292730 219218 292966 219454
rect 292730 218898 292966 219134
rect 293546 186618 294102 187174
rect 289826 182898 290382 183454
rect 292730 183218 292966 183454
rect 292730 182898 292966 183134
rect 293546 150618 294102 151174
rect 289826 146898 290382 147454
rect 292730 147218 292966 147454
rect 292730 146898 292966 147134
rect 293546 114618 294102 115174
rect 289826 110898 290382 111454
rect 292730 111218 292966 111454
rect 292730 110898 292966 111134
rect 293546 78618 294102 79174
rect 289826 74898 290382 75454
rect 292730 75218 292966 75454
rect 292730 74898 292966 75134
rect 293546 42618 294102 43174
rect 289826 38898 290382 39454
rect 292730 39218 292966 39454
rect 292730 38898 292966 39134
rect 289826 2898 290382 3454
rect 289826 -902 290382 -346
rect 293546 6618 294102 7174
rect 293546 -1862 294102 -1306
rect 297266 706202 297822 706758
rect 297266 694338 297822 694894
rect 297266 658338 297822 658894
rect 297266 622338 297822 622894
rect 297266 586338 297822 586894
rect 297266 550338 297822 550894
rect 297266 514338 297822 514894
rect 297266 478338 297822 478894
rect 297266 442338 297822 442894
rect 297266 406338 297822 406894
rect 297266 370338 297822 370894
rect 297266 334338 297822 334894
rect 297266 298338 297822 298894
rect 297266 262338 297822 262894
rect 297266 226338 297822 226894
rect 297266 190338 297822 190894
rect 297266 154338 297822 154894
rect 297266 118338 297822 118894
rect 297266 82338 297822 82894
rect 297266 46338 297822 46894
rect 297266 10338 297822 10894
rect 297266 -2822 297822 -2266
rect 300986 707162 301542 707718
rect 300986 698058 301542 698614
rect 300986 662058 301542 662614
rect 300986 626058 301542 626614
rect 300986 590058 301542 590614
rect 300986 554058 301542 554614
rect 300986 518058 301542 518614
rect 300986 482058 301542 482614
rect 300986 446058 301542 446614
rect 300986 410058 301542 410614
rect 300986 374058 301542 374614
rect 300986 338058 301542 338614
rect 300986 302058 301542 302614
rect 300986 266058 301542 266614
rect 300986 230058 301542 230614
rect 300986 194058 301542 194614
rect 300986 158058 301542 158614
rect 300986 122058 301542 122614
rect 300986 86058 301542 86614
rect 300986 50058 301542 50614
rect 300986 14058 301542 14614
rect 300986 -3782 301542 -3226
rect 304706 708122 305262 708678
rect 304706 665778 305262 666334
rect 304706 629778 305262 630334
rect 304706 593778 305262 594334
rect 304706 557778 305262 558334
rect 304706 521778 305262 522334
rect 304706 485778 305262 486334
rect 304706 449778 305262 450334
rect 304706 413778 305262 414334
rect 304706 377778 305262 378334
rect 308426 709082 308982 709638
rect 308426 669498 308982 670054
rect 308426 633498 308982 634054
rect 308426 597498 308982 598054
rect 308426 561498 308982 562054
rect 308426 525498 308982 526054
rect 308426 489498 308982 490054
rect 308426 453498 308982 454054
rect 308426 417498 308982 418054
rect 308426 381498 308982 382054
rect 312146 710042 312702 710598
rect 312146 673218 312702 673774
rect 312146 637218 312702 637774
rect 312146 601218 312702 601774
rect 312146 565218 312702 565774
rect 312146 529218 312702 529774
rect 312146 493218 312702 493774
rect 312146 457218 312702 457774
rect 312146 421218 312702 421774
rect 312146 385218 312702 385774
rect 304706 341778 305262 342334
rect 312146 349218 312702 349774
rect 308090 330938 308326 331174
rect 308090 330618 308326 330854
rect 304706 305778 305262 306334
rect 312146 313218 312702 313774
rect 308090 294938 308326 295174
rect 308090 294618 308326 294854
rect 304706 269778 305262 270334
rect 312146 277218 312702 277774
rect 308090 258938 308326 259174
rect 308090 258618 308326 258854
rect 304706 233778 305262 234334
rect 312146 241218 312702 241774
rect 308090 222938 308326 223174
rect 308090 222618 308326 222854
rect 304706 197778 305262 198334
rect 312146 205218 312702 205774
rect 308090 186938 308326 187174
rect 308090 186618 308326 186854
rect 304706 161778 305262 162334
rect 312146 169218 312702 169774
rect 308090 150938 308326 151174
rect 308090 150618 308326 150854
rect 304706 125778 305262 126334
rect 312146 133218 312702 133774
rect 308090 114938 308326 115174
rect 308090 114618 308326 114854
rect 304706 89778 305262 90334
rect 312146 97218 312702 97774
rect 308090 78938 308326 79174
rect 308090 78618 308326 78854
rect 304706 53778 305262 54334
rect 312146 61218 312702 61774
rect 308090 42938 308326 43174
rect 308090 42618 308326 42854
rect 304706 17778 305262 18334
rect 312146 25218 312702 25774
rect 308090 6938 308326 7174
rect 308090 6618 308326 6854
rect 304706 -4742 305262 -4186
rect 312146 -6662 312702 -6106
rect 315866 711002 316422 711558
rect 315866 676938 316422 677494
rect 315866 640938 316422 641494
rect 315866 604938 316422 605494
rect 315866 568938 316422 569494
rect 315866 532938 316422 533494
rect 315866 496938 316422 497494
rect 315866 460938 316422 461494
rect 315866 424938 316422 425494
rect 315866 388938 316422 389494
rect 315866 352938 316422 353494
rect 325826 704282 326382 704838
rect 325826 686898 326382 687454
rect 325826 650898 326382 651454
rect 325826 614898 326382 615454
rect 325826 578898 326382 579454
rect 325826 542898 326382 543454
rect 325826 506898 326382 507454
rect 325826 470898 326382 471454
rect 325826 434898 326382 435454
rect 325826 398898 326382 399454
rect 325826 362898 326382 363454
rect 323450 327218 323686 327454
rect 323450 326898 323686 327134
rect 325826 326898 326382 327454
rect 315866 316938 316422 317494
rect 323450 291218 323686 291454
rect 323450 290898 323686 291134
rect 325826 290898 326382 291454
rect 315866 280938 316422 281494
rect 323450 255218 323686 255454
rect 323450 254898 323686 255134
rect 325826 254898 326382 255454
rect 315866 244938 316422 245494
rect 323450 219218 323686 219454
rect 323450 218898 323686 219134
rect 325826 218898 326382 219454
rect 315866 208938 316422 209494
rect 323450 183218 323686 183454
rect 323450 182898 323686 183134
rect 325826 182898 326382 183454
rect 315866 172938 316422 173494
rect 323450 147218 323686 147454
rect 323450 146898 323686 147134
rect 325826 146898 326382 147454
rect 315866 136938 316422 137494
rect 323450 111218 323686 111454
rect 323450 110898 323686 111134
rect 325826 110898 326382 111454
rect 315866 100938 316422 101494
rect 323450 75218 323686 75454
rect 323450 74898 323686 75134
rect 325826 74898 326382 75454
rect 315866 64938 316422 65494
rect 323450 39218 323686 39454
rect 323450 38898 323686 39134
rect 325826 38898 326382 39454
rect 315866 28938 316422 29494
rect 315866 -7622 316422 -7066
rect 325826 2898 326382 3454
rect 325826 -902 326382 -346
rect 329546 705242 330102 705798
rect 329546 690618 330102 691174
rect 329546 654618 330102 655174
rect 329546 618618 330102 619174
rect 329546 582618 330102 583174
rect 329546 546618 330102 547174
rect 329546 510618 330102 511174
rect 329546 474618 330102 475174
rect 329546 438618 330102 439174
rect 329546 402618 330102 403174
rect 329546 366618 330102 367174
rect 329546 330618 330102 331174
rect 329546 294618 330102 295174
rect 329546 258618 330102 259174
rect 329546 222618 330102 223174
rect 329546 186618 330102 187174
rect 329546 150618 330102 151174
rect 329546 114618 330102 115174
rect 329546 78618 330102 79174
rect 329546 42618 330102 43174
rect 329546 6618 330102 7174
rect 329546 -1862 330102 -1306
rect 333266 706202 333822 706758
rect 333266 694338 333822 694894
rect 333266 658338 333822 658894
rect 333266 622338 333822 622894
rect 333266 586338 333822 586894
rect 333266 550338 333822 550894
rect 333266 514338 333822 514894
rect 333266 478338 333822 478894
rect 333266 442338 333822 442894
rect 333266 406338 333822 406894
rect 333266 370338 333822 370894
rect 333266 334338 333822 334894
rect 333266 298338 333822 298894
rect 333266 262338 333822 262894
rect 333266 226338 333822 226894
rect 333266 190338 333822 190894
rect 333266 154338 333822 154894
rect 333266 118338 333822 118894
rect 333266 82338 333822 82894
rect 333266 46338 333822 46894
rect 333266 10338 333822 10894
rect 333266 -2822 333822 -2266
rect 336986 707162 337542 707718
rect 336986 698058 337542 698614
rect 336986 662058 337542 662614
rect 336986 626058 337542 626614
rect 336986 590058 337542 590614
rect 336986 554058 337542 554614
rect 336986 518058 337542 518614
rect 336986 482058 337542 482614
rect 336986 446058 337542 446614
rect 336986 410058 337542 410614
rect 336986 374058 337542 374614
rect 336986 338058 337542 338614
rect 340706 708122 341262 708678
rect 340706 665778 341262 666334
rect 340706 629778 341262 630334
rect 340706 593778 341262 594334
rect 340706 557778 341262 558334
rect 340706 521778 341262 522334
rect 340706 485778 341262 486334
rect 340706 449778 341262 450334
rect 340706 413778 341262 414334
rect 340706 377778 341262 378334
rect 340706 341778 341262 342334
rect 338810 330938 339046 331174
rect 338810 330618 339046 330854
rect 336986 302058 337542 302614
rect 340706 305778 341262 306334
rect 338810 294938 339046 295174
rect 338810 294618 339046 294854
rect 336986 266058 337542 266614
rect 340706 269778 341262 270334
rect 338810 258938 339046 259174
rect 338810 258618 339046 258854
rect 336986 230058 337542 230614
rect 340706 233778 341262 234334
rect 338810 222938 339046 223174
rect 338810 222618 339046 222854
rect 336986 194058 337542 194614
rect 340706 197778 341262 198334
rect 338810 186938 339046 187174
rect 338810 186618 339046 186854
rect 336986 158058 337542 158614
rect 340706 161778 341262 162334
rect 338810 150938 339046 151174
rect 338810 150618 339046 150854
rect 336986 122058 337542 122614
rect 340706 125778 341262 126334
rect 338810 114938 339046 115174
rect 338810 114618 339046 114854
rect 336986 86058 337542 86614
rect 340706 89778 341262 90334
rect 338810 78938 339046 79174
rect 338810 78618 339046 78854
rect 336986 50058 337542 50614
rect 340706 53778 341262 54334
rect 338810 42938 339046 43174
rect 338810 42618 339046 42854
rect 336986 14058 337542 14614
rect 340706 17778 341262 18334
rect 338810 6938 339046 7174
rect 338810 6618 339046 6854
rect 336986 -3782 337542 -3226
rect 340706 -4742 341262 -4186
rect 344426 709082 344982 709638
rect 344426 669498 344982 670054
rect 344426 633498 344982 634054
rect 344426 597498 344982 598054
rect 344426 561498 344982 562054
rect 344426 525498 344982 526054
rect 344426 489498 344982 490054
rect 344426 453498 344982 454054
rect 344426 417498 344982 418054
rect 344426 381498 344982 382054
rect 344426 345498 344982 346054
rect 344426 309498 344982 310054
rect 344426 273498 344982 274054
rect 344426 237498 344982 238054
rect 344426 201498 344982 202054
rect 344426 165498 344982 166054
rect 344426 129498 344982 130054
rect 344426 93498 344982 94054
rect 344426 57498 344982 58054
rect 344426 21498 344982 22054
rect 344426 -5702 344982 -5146
rect 348146 710042 348702 710598
rect 348146 673218 348702 673774
rect 348146 637218 348702 637774
rect 348146 601218 348702 601774
rect 348146 565218 348702 565774
rect 348146 529218 348702 529774
rect 348146 493218 348702 493774
rect 348146 457218 348702 457774
rect 348146 421218 348702 421774
rect 348146 385218 348702 385774
rect 348146 349218 348702 349774
rect 348146 313218 348702 313774
rect 348146 277218 348702 277774
rect 348146 241218 348702 241774
rect 348146 205218 348702 205774
rect 348146 169218 348702 169774
rect 348146 133218 348702 133774
rect 348146 97218 348702 97774
rect 348146 61218 348702 61774
rect 348146 25218 348702 25774
rect 348146 -6662 348702 -6106
rect 351866 711002 352422 711558
rect 351866 676938 352422 677494
rect 351866 640938 352422 641494
rect 351866 604938 352422 605494
rect 351866 568938 352422 569494
rect 351866 532938 352422 533494
rect 351866 496938 352422 497494
rect 351866 460938 352422 461494
rect 351866 424938 352422 425494
rect 351866 388938 352422 389494
rect 351866 352938 352422 353494
rect 361826 704282 362382 704838
rect 361826 686898 362382 687454
rect 361826 650898 362382 651454
rect 361826 614898 362382 615454
rect 361826 578898 362382 579454
rect 361826 542898 362382 543454
rect 361826 506898 362382 507454
rect 361826 470898 362382 471454
rect 361826 434898 362382 435454
rect 361826 398898 362382 399454
rect 361826 362898 362382 363454
rect 354170 327218 354406 327454
rect 354170 326898 354406 327134
rect 361826 326898 362382 327454
rect 351866 316938 352422 317494
rect 354170 291218 354406 291454
rect 354170 290898 354406 291134
rect 361826 290898 362382 291454
rect 351866 280938 352422 281494
rect 354170 255218 354406 255454
rect 354170 254898 354406 255134
rect 361826 254898 362382 255454
rect 351866 244938 352422 245494
rect 354170 219218 354406 219454
rect 354170 218898 354406 219134
rect 361826 218898 362382 219454
rect 351866 208938 352422 209494
rect 354170 183218 354406 183454
rect 354170 182898 354406 183134
rect 361826 182898 362382 183454
rect 351866 172938 352422 173494
rect 354170 147218 354406 147454
rect 354170 146898 354406 147134
rect 361826 146898 362382 147454
rect 351866 136938 352422 137494
rect 354170 111218 354406 111454
rect 354170 110898 354406 111134
rect 361826 110898 362382 111454
rect 351866 100938 352422 101494
rect 354170 75218 354406 75454
rect 354170 74898 354406 75134
rect 361826 74898 362382 75454
rect 351866 64938 352422 65494
rect 354170 39218 354406 39454
rect 354170 38898 354406 39134
rect 361826 38898 362382 39454
rect 351866 28938 352422 29494
rect 351866 -7622 352422 -7066
rect 361826 2898 362382 3454
rect 365546 705242 366102 705798
rect 365546 690618 366102 691174
rect 365546 654618 366102 655174
rect 365546 618618 366102 619174
rect 365546 582618 366102 583174
rect 365546 546618 366102 547174
rect 365546 510618 366102 511174
rect 365546 474618 366102 475174
rect 365546 438618 366102 439174
rect 365546 402618 366102 403174
rect 365546 366618 366102 367174
rect 369266 706202 369822 706758
rect 369266 694338 369822 694894
rect 369266 658338 369822 658894
rect 369266 622338 369822 622894
rect 369266 586338 369822 586894
rect 369266 550338 369822 550894
rect 369266 514338 369822 514894
rect 369266 478338 369822 478894
rect 369266 442338 369822 442894
rect 369266 406338 369822 406894
rect 369266 370338 369822 370894
rect 372986 707162 373542 707718
rect 372986 698058 373542 698614
rect 372986 662058 373542 662614
rect 372986 626058 373542 626614
rect 372986 590058 373542 590614
rect 372986 554058 373542 554614
rect 372986 518058 373542 518614
rect 372986 482058 373542 482614
rect 372986 446058 373542 446614
rect 372986 410058 373542 410614
rect 372986 374058 373542 374614
rect 372986 338058 373542 338614
rect 365546 330618 366102 331174
rect 369530 330938 369766 331174
rect 369530 330618 369766 330854
rect 372986 302058 373542 302614
rect 365546 294618 366102 295174
rect 369530 294938 369766 295174
rect 369530 294618 369766 294854
rect 372986 266058 373542 266614
rect 365546 258618 366102 259174
rect 369530 258938 369766 259174
rect 369530 258618 369766 258854
rect 372986 230058 373542 230614
rect 365546 222618 366102 223174
rect 369530 222938 369766 223174
rect 369530 222618 369766 222854
rect 372986 194058 373542 194614
rect 365546 186618 366102 187174
rect 369530 186938 369766 187174
rect 369530 186618 369766 186854
rect 372986 158058 373542 158614
rect 365546 150618 366102 151174
rect 369530 150938 369766 151174
rect 369530 150618 369766 150854
rect 372986 122058 373542 122614
rect 365546 114618 366102 115174
rect 369530 114938 369766 115174
rect 369530 114618 369766 114854
rect 372986 86058 373542 86614
rect 365546 78618 366102 79174
rect 369530 78938 369766 79174
rect 369530 78618 369766 78854
rect 372986 50058 373542 50614
rect 365546 42618 366102 43174
rect 369530 42938 369766 43174
rect 369530 42618 369766 42854
rect 372986 14058 373542 14614
rect 365546 6618 366102 7174
rect 361826 -902 362382 -346
rect 369530 6938 369766 7174
rect 369530 6618 369766 6854
rect 365546 -1862 366102 -1306
rect 372986 -3782 373542 -3226
rect 376706 708122 377262 708678
rect 376706 665778 377262 666334
rect 376706 629778 377262 630334
rect 376706 593778 377262 594334
rect 376706 557778 377262 558334
rect 376706 521778 377262 522334
rect 376706 485778 377262 486334
rect 376706 449778 377262 450334
rect 376706 413778 377262 414334
rect 376706 377778 377262 378334
rect 376706 341778 377262 342334
rect 376706 305778 377262 306334
rect 376706 269778 377262 270334
rect 376706 233778 377262 234334
rect 376706 197778 377262 198334
rect 376706 161778 377262 162334
rect 376706 125778 377262 126334
rect 376706 89778 377262 90334
rect 376706 53778 377262 54334
rect 376706 17778 377262 18334
rect 380426 709082 380982 709638
rect 380426 669498 380982 670054
rect 380426 633498 380982 634054
rect 380426 597498 380982 598054
rect 380426 561498 380982 562054
rect 380426 525498 380982 526054
rect 380426 489498 380982 490054
rect 380426 453498 380982 454054
rect 380426 417498 380982 418054
rect 380426 381498 380982 382054
rect 384146 710042 384702 710598
rect 384146 673218 384702 673774
rect 384146 637218 384702 637774
rect 384146 601218 384702 601774
rect 384146 565218 384702 565774
rect 384146 529218 384702 529774
rect 384146 493218 384702 493774
rect 384146 457218 384702 457774
rect 384146 421218 384702 421774
rect 384146 385218 384702 385774
rect 387866 711002 388422 711558
rect 387866 676938 388422 677494
rect 387866 640938 388422 641494
rect 387866 604938 388422 605494
rect 387866 568938 388422 569494
rect 387866 532938 388422 533494
rect 387866 496938 388422 497494
rect 387866 460938 388422 461494
rect 387866 424938 388422 425494
rect 387866 388938 388422 389494
rect 380426 345498 380982 346054
rect 387866 352938 388422 353494
rect 384890 327218 385126 327454
rect 384890 326898 385126 327134
rect 380426 309498 380982 310054
rect 387866 316938 388422 317494
rect 384890 291218 385126 291454
rect 384890 290898 385126 291134
rect 380426 273498 380982 274054
rect 387866 280938 388422 281494
rect 384890 255218 385126 255454
rect 384890 254898 385126 255134
rect 380426 237498 380982 238054
rect 387866 244938 388422 245494
rect 384890 219218 385126 219454
rect 384890 218898 385126 219134
rect 380426 201498 380982 202054
rect 387866 208938 388422 209494
rect 384890 183218 385126 183454
rect 384890 182898 385126 183134
rect 380426 165498 380982 166054
rect 387866 172938 388422 173494
rect 384890 147218 385126 147454
rect 384890 146898 385126 147134
rect 380426 129498 380982 130054
rect 387866 136938 388422 137494
rect 384890 111218 385126 111454
rect 384890 110898 385126 111134
rect 380426 93498 380982 94054
rect 387866 100938 388422 101494
rect 384890 75218 385126 75454
rect 384890 74898 385126 75134
rect 380426 57498 380982 58054
rect 387866 64938 388422 65494
rect 384890 39218 385126 39454
rect 384890 38898 385126 39134
rect 380426 21498 380982 22054
rect 376706 -4742 377262 -4186
rect 387866 28938 388422 29494
rect 380426 -5702 380982 -5146
rect 397826 704282 398382 704838
rect 397826 686898 398382 687454
rect 397826 650898 398382 651454
rect 397826 614898 398382 615454
rect 397826 578898 398382 579454
rect 397826 542898 398382 543454
rect 397826 506898 398382 507454
rect 397826 470898 398382 471454
rect 397826 434898 398382 435454
rect 397826 398898 398382 399454
rect 397826 362898 398382 363454
rect 401546 705242 402102 705798
rect 401546 690618 402102 691174
rect 401546 654618 402102 655174
rect 401546 618618 402102 619174
rect 401546 582618 402102 583174
rect 401546 546618 402102 547174
rect 401546 510618 402102 511174
rect 401546 474618 402102 475174
rect 401546 438618 402102 439174
rect 401546 402618 402102 403174
rect 401546 366618 402102 367174
rect 400250 330938 400486 331174
rect 400250 330618 400486 330854
rect 401546 330618 402102 331174
rect 397826 326898 398382 327454
rect 400250 294938 400486 295174
rect 400250 294618 400486 294854
rect 401546 294618 402102 295174
rect 397826 290898 398382 291454
rect 400250 258938 400486 259174
rect 400250 258618 400486 258854
rect 401546 258618 402102 259174
rect 397826 254898 398382 255454
rect 400250 222938 400486 223174
rect 400250 222618 400486 222854
rect 401546 222618 402102 223174
rect 397826 218898 398382 219454
rect 400250 186938 400486 187174
rect 400250 186618 400486 186854
rect 401546 186618 402102 187174
rect 397826 182898 398382 183454
rect 400250 150938 400486 151174
rect 400250 150618 400486 150854
rect 401546 150618 402102 151174
rect 397826 146898 398382 147454
rect 400250 114938 400486 115174
rect 400250 114618 400486 114854
rect 401546 114618 402102 115174
rect 397826 110898 398382 111454
rect 400250 78938 400486 79174
rect 400250 78618 400486 78854
rect 401546 78618 402102 79174
rect 397826 74898 398382 75454
rect 400250 42938 400486 43174
rect 400250 42618 400486 42854
rect 401546 42618 402102 43174
rect 397826 38898 398382 39454
rect 400250 6938 400486 7174
rect 400250 6618 400486 6854
rect 401546 6618 402102 7174
rect 397826 2898 398382 3454
rect 387866 -7622 388422 -7066
rect 397826 -902 398382 -346
rect 401546 -1862 402102 -1306
rect 405266 706202 405822 706758
rect 405266 694338 405822 694894
rect 405266 658338 405822 658894
rect 405266 622338 405822 622894
rect 405266 586338 405822 586894
rect 405266 550338 405822 550894
rect 405266 514338 405822 514894
rect 405266 478338 405822 478894
rect 405266 442338 405822 442894
rect 405266 406338 405822 406894
rect 405266 370338 405822 370894
rect 405266 334338 405822 334894
rect 405266 298338 405822 298894
rect 405266 262338 405822 262894
rect 405266 226338 405822 226894
rect 405266 190338 405822 190894
rect 405266 154338 405822 154894
rect 405266 118338 405822 118894
rect 405266 82338 405822 82894
rect 405266 46338 405822 46894
rect 405266 10338 405822 10894
rect 408986 707162 409542 707718
rect 408986 698058 409542 698614
rect 408986 662058 409542 662614
rect 408986 626058 409542 626614
rect 408986 590058 409542 590614
rect 408986 554058 409542 554614
rect 408986 518058 409542 518614
rect 408986 482058 409542 482614
rect 408986 446058 409542 446614
rect 408986 410058 409542 410614
rect 408986 374058 409542 374614
rect 408986 338058 409542 338614
rect 408986 302058 409542 302614
rect 408986 266058 409542 266614
rect 408986 230058 409542 230614
rect 408986 194058 409542 194614
rect 408986 158058 409542 158614
rect 408986 122058 409542 122614
rect 408986 86058 409542 86614
rect 408986 50058 409542 50614
rect 408986 14058 409542 14614
rect 405266 -2822 405822 -2266
rect 408986 -3782 409542 -3226
rect 412706 708122 413262 708678
rect 412706 665778 413262 666334
rect 412706 629778 413262 630334
rect 412706 593778 413262 594334
rect 412706 557778 413262 558334
rect 412706 521778 413262 522334
rect 412706 485778 413262 486334
rect 412706 449778 413262 450334
rect 412706 413778 413262 414334
rect 412706 377778 413262 378334
rect 412706 341778 413262 342334
rect 416426 709082 416982 709638
rect 416426 669498 416982 670054
rect 416426 633498 416982 634054
rect 416426 597498 416982 598054
rect 416426 561498 416982 562054
rect 416426 525498 416982 526054
rect 416426 489498 416982 490054
rect 416426 453498 416982 454054
rect 416426 417498 416982 418054
rect 416426 381498 416982 382054
rect 416426 345498 416982 346054
rect 415610 327218 415846 327454
rect 415610 326898 415846 327134
rect 412706 305778 413262 306334
rect 416426 309498 416982 310054
rect 415610 291218 415846 291454
rect 415610 290898 415846 291134
rect 412706 269778 413262 270334
rect 416426 273498 416982 274054
rect 415610 255218 415846 255454
rect 415610 254898 415846 255134
rect 412706 233778 413262 234334
rect 416426 237498 416982 238054
rect 415610 219218 415846 219454
rect 415610 218898 415846 219134
rect 412706 197778 413262 198334
rect 416426 201498 416982 202054
rect 415610 183218 415846 183454
rect 415610 182898 415846 183134
rect 412706 161778 413262 162334
rect 416426 165498 416982 166054
rect 415610 147218 415846 147454
rect 415610 146898 415846 147134
rect 412706 125778 413262 126334
rect 416426 129498 416982 130054
rect 415610 111218 415846 111454
rect 415610 110898 415846 111134
rect 412706 89778 413262 90334
rect 416426 93498 416982 94054
rect 415610 75218 415846 75454
rect 415610 74898 415846 75134
rect 412706 53778 413262 54334
rect 416426 57498 416982 58054
rect 415610 39218 415846 39454
rect 415610 38898 415846 39134
rect 412706 17778 413262 18334
rect 412706 -4742 413262 -4186
rect 416426 21498 416982 22054
rect 416426 -5702 416982 -5146
rect 420146 710042 420702 710598
rect 420146 673218 420702 673774
rect 420146 637218 420702 637774
rect 420146 601218 420702 601774
rect 420146 565218 420702 565774
rect 420146 529218 420702 529774
rect 420146 493218 420702 493774
rect 420146 457218 420702 457774
rect 420146 421218 420702 421774
rect 420146 385218 420702 385774
rect 420146 349218 420702 349774
rect 420146 313218 420702 313774
rect 420146 277218 420702 277774
rect 420146 241218 420702 241774
rect 420146 205218 420702 205774
rect 420146 169218 420702 169774
rect 420146 133218 420702 133774
rect 420146 97218 420702 97774
rect 420146 61218 420702 61774
rect 420146 25218 420702 25774
rect 420146 -6662 420702 -6106
rect 423866 711002 424422 711558
rect 423866 676938 424422 677494
rect 423866 640938 424422 641494
rect 423866 604938 424422 605494
rect 423866 568938 424422 569494
rect 423866 532938 424422 533494
rect 423866 496938 424422 497494
rect 423866 460938 424422 461494
rect 423866 424938 424422 425494
rect 423866 388938 424422 389494
rect 423866 352938 424422 353494
rect 433826 704282 434382 704838
rect 433826 686898 434382 687454
rect 433826 650898 434382 651454
rect 433826 614898 434382 615454
rect 433826 578898 434382 579454
rect 433826 542898 434382 543454
rect 433826 506898 434382 507454
rect 433826 470898 434382 471454
rect 433826 434898 434382 435454
rect 433826 398898 434382 399454
rect 433826 362898 434382 363454
rect 430970 330938 431206 331174
rect 430970 330618 431206 330854
rect 423866 316938 424422 317494
rect 433826 326898 434382 327454
rect 430970 294938 431206 295174
rect 430970 294618 431206 294854
rect 423866 280938 424422 281494
rect 433826 290898 434382 291454
rect 430970 258938 431206 259174
rect 430970 258618 431206 258854
rect 423866 244938 424422 245494
rect 433826 254898 434382 255454
rect 430970 222938 431206 223174
rect 430970 222618 431206 222854
rect 423866 208938 424422 209494
rect 433826 218898 434382 219454
rect 430970 186938 431206 187174
rect 430970 186618 431206 186854
rect 423866 172938 424422 173494
rect 433826 182898 434382 183454
rect 430970 150938 431206 151174
rect 430970 150618 431206 150854
rect 423866 136938 424422 137494
rect 433826 146898 434382 147454
rect 430970 114938 431206 115174
rect 430970 114618 431206 114854
rect 423866 100938 424422 101494
rect 433826 110898 434382 111454
rect 430970 78938 431206 79174
rect 430970 78618 431206 78854
rect 423866 64938 424422 65494
rect 433826 74898 434382 75454
rect 430970 42938 431206 43174
rect 430970 42618 431206 42854
rect 423866 28938 424422 29494
rect 433826 38898 434382 39454
rect 430970 6938 431206 7174
rect 430970 6618 431206 6854
rect 423866 -7622 424422 -7066
rect 433826 2898 434382 3454
rect 433826 -902 434382 -346
rect 437546 705242 438102 705798
rect 437546 690618 438102 691174
rect 437546 654618 438102 655174
rect 437546 618618 438102 619174
rect 437546 582618 438102 583174
rect 437546 546618 438102 547174
rect 437546 510618 438102 511174
rect 437546 474618 438102 475174
rect 437546 438618 438102 439174
rect 437546 402618 438102 403174
rect 437546 366618 438102 367174
rect 437546 330618 438102 331174
rect 437546 294618 438102 295174
rect 437546 258618 438102 259174
rect 437546 222618 438102 223174
rect 437546 186618 438102 187174
rect 437546 150618 438102 151174
rect 437546 114618 438102 115174
rect 437546 78618 438102 79174
rect 437546 42618 438102 43174
rect 437546 6618 438102 7174
rect 437546 -1862 438102 -1306
rect 441266 706202 441822 706758
rect 441266 694338 441822 694894
rect 441266 658338 441822 658894
rect 441266 622338 441822 622894
rect 441266 586338 441822 586894
rect 441266 550338 441822 550894
rect 441266 514338 441822 514894
rect 441266 478338 441822 478894
rect 441266 442338 441822 442894
rect 441266 406338 441822 406894
rect 441266 370338 441822 370894
rect 441266 334338 441822 334894
rect 441266 298338 441822 298894
rect 441266 262338 441822 262894
rect 441266 226338 441822 226894
rect 441266 190338 441822 190894
rect 441266 154338 441822 154894
rect 441266 118338 441822 118894
rect 441266 82338 441822 82894
rect 441266 46338 441822 46894
rect 441266 10338 441822 10894
rect 441266 -2822 441822 -2266
rect 444986 707162 445542 707718
rect 444986 698058 445542 698614
rect 444986 662058 445542 662614
rect 444986 626058 445542 626614
rect 444986 590058 445542 590614
rect 444986 554058 445542 554614
rect 444986 518058 445542 518614
rect 444986 482058 445542 482614
rect 444986 446058 445542 446614
rect 444986 410058 445542 410614
rect 444986 374058 445542 374614
rect 444986 338058 445542 338614
rect 448706 708122 449262 708678
rect 448706 665778 449262 666334
rect 448706 629778 449262 630334
rect 448706 593778 449262 594334
rect 448706 557778 449262 558334
rect 448706 521778 449262 522334
rect 448706 485778 449262 486334
rect 448706 449778 449262 450334
rect 448706 413778 449262 414334
rect 448706 377778 449262 378334
rect 448706 341778 449262 342334
rect 446330 327218 446566 327454
rect 446330 326898 446566 327134
rect 444986 302058 445542 302614
rect 448706 305778 449262 306334
rect 446330 291218 446566 291454
rect 446330 290898 446566 291134
rect 444986 266058 445542 266614
rect 448706 269778 449262 270334
rect 446330 255218 446566 255454
rect 446330 254898 446566 255134
rect 444986 230058 445542 230614
rect 448706 233778 449262 234334
rect 446330 219218 446566 219454
rect 446330 218898 446566 219134
rect 444986 194058 445542 194614
rect 448706 197778 449262 198334
rect 446330 183218 446566 183454
rect 446330 182898 446566 183134
rect 444986 158058 445542 158614
rect 448706 161778 449262 162334
rect 446330 147218 446566 147454
rect 446330 146898 446566 147134
rect 444986 122058 445542 122614
rect 448706 125778 449262 126334
rect 446330 111218 446566 111454
rect 446330 110898 446566 111134
rect 444986 86058 445542 86614
rect 448706 89778 449262 90334
rect 446330 75218 446566 75454
rect 446330 74898 446566 75134
rect 444986 50058 445542 50614
rect 448706 53778 449262 54334
rect 446330 39218 446566 39454
rect 446330 38898 446566 39134
rect 444986 14058 445542 14614
rect 444986 -3782 445542 -3226
rect 448706 17778 449262 18334
rect 448706 -4742 449262 -4186
rect 452426 709082 452982 709638
rect 452426 669498 452982 670054
rect 452426 633498 452982 634054
rect 452426 597498 452982 598054
rect 452426 561498 452982 562054
rect 452426 525498 452982 526054
rect 452426 489498 452982 490054
rect 452426 453498 452982 454054
rect 452426 417498 452982 418054
rect 452426 381498 452982 382054
rect 452426 345498 452982 346054
rect 452426 309498 452982 310054
rect 452426 273498 452982 274054
rect 452426 237498 452982 238054
rect 452426 201498 452982 202054
rect 452426 165498 452982 166054
rect 452426 129498 452982 130054
rect 452426 93498 452982 94054
rect 452426 57498 452982 58054
rect 452426 21498 452982 22054
rect 452426 -5702 452982 -5146
rect 456146 710042 456702 710598
rect 456146 673218 456702 673774
rect 456146 637218 456702 637774
rect 456146 601218 456702 601774
rect 456146 565218 456702 565774
rect 456146 529218 456702 529774
rect 456146 493218 456702 493774
rect 456146 457218 456702 457774
rect 456146 421218 456702 421774
rect 456146 385218 456702 385774
rect 456146 349218 456702 349774
rect 456146 313218 456702 313774
rect 456146 277218 456702 277774
rect 456146 241218 456702 241774
rect 456146 205218 456702 205774
rect 456146 169218 456702 169774
rect 456146 133218 456702 133774
rect 456146 97218 456702 97774
rect 456146 61218 456702 61774
rect 456146 25218 456702 25774
rect 459866 711002 460422 711558
rect 459866 676938 460422 677494
rect 459866 640938 460422 641494
rect 459866 604938 460422 605494
rect 459866 568938 460422 569494
rect 459866 532938 460422 533494
rect 459866 496938 460422 497494
rect 459866 460938 460422 461494
rect 459866 424938 460422 425494
rect 459866 388938 460422 389494
rect 459866 352938 460422 353494
rect 469826 704282 470382 704838
rect 469826 686898 470382 687454
rect 469826 650898 470382 651454
rect 469826 614898 470382 615454
rect 469826 578898 470382 579454
rect 469826 542898 470382 543454
rect 469826 506898 470382 507454
rect 469826 470898 470382 471454
rect 469826 434898 470382 435454
rect 469826 398898 470382 399454
rect 469826 362898 470382 363454
rect 461690 330938 461926 331174
rect 461690 330618 461926 330854
rect 459866 316938 460422 317494
rect 469826 326898 470382 327454
rect 461690 294938 461926 295174
rect 461690 294618 461926 294854
rect 459866 280938 460422 281494
rect 469826 290898 470382 291454
rect 461690 258938 461926 259174
rect 461690 258618 461926 258854
rect 459866 244938 460422 245494
rect 469826 254898 470382 255454
rect 461690 222938 461926 223174
rect 461690 222618 461926 222854
rect 459866 208938 460422 209494
rect 469826 218898 470382 219454
rect 461690 186938 461926 187174
rect 461690 186618 461926 186854
rect 459866 172938 460422 173494
rect 469826 182898 470382 183454
rect 461690 150938 461926 151174
rect 461690 150618 461926 150854
rect 459866 136938 460422 137494
rect 469826 146898 470382 147454
rect 461690 114938 461926 115174
rect 461690 114618 461926 114854
rect 459866 100938 460422 101494
rect 469826 110898 470382 111454
rect 461690 78938 461926 79174
rect 461690 78618 461926 78854
rect 459866 64938 460422 65494
rect 469826 74898 470382 75454
rect 461690 42938 461926 43174
rect 461690 42618 461926 42854
rect 459866 28938 460422 29494
rect 456146 -6662 456702 -6106
rect 469826 38898 470382 39454
rect 461690 6938 461926 7174
rect 461690 6618 461926 6854
rect 469826 2898 470382 3454
rect 459866 -7622 460422 -7066
rect 469826 -902 470382 -346
rect 473546 705242 474102 705798
rect 473546 690618 474102 691174
rect 473546 654618 474102 655174
rect 473546 618618 474102 619174
rect 473546 582618 474102 583174
rect 473546 546618 474102 547174
rect 473546 510618 474102 511174
rect 473546 474618 474102 475174
rect 473546 438618 474102 439174
rect 473546 402618 474102 403174
rect 473546 366618 474102 367174
rect 477266 706202 477822 706758
rect 477266 694338 477822 694894
rect 477266 658338 477822 658894
rect 477266 622338 477822 622894
rect 477266 586338 477822 586894
rect 477266 550338 477822 550894
rect 477266 514338 477822 514894
rect 477266 478338 477822 478894
rect 477266 442338 477822 442894
rect 477266 406338 477822 406894
rect 477266 370338 477822 370894
rect 480986 707162 481542 707718
rect 480986 698058 481542 698614
rect 480986 662058 481542 662614
rect 480986 626058 481542 626614
rect 480986 590058 481542 590614
rect 480986 554058 481542 554614
rect 480986 518058 481542 518614
rect 480986 482058 481542 482614
rect 480986 446058 481542 446614
rect 480986 410058 481542 410614
rect 480986 374058 481542 374614
rect 473546 330618 474102 331174
rect 480986 338058 481542 338614
rect 477050 327218 477286 327454
rect 477050 326898 477286 327134
rect 473546 294618 474102 295174
rect 480986 302058 481542 302614
rect 477050 291218 477286 291454
rect 477050 290898 477286 291134
rect 473546 258618 474102 259174
rect 480986 266058 481542 266614
rect 477050 255218 477286 255454
rect 477050 254898 477286 255134
rect 473546 222618 474102 223174
rect 480986 230058 481542 230614
rect 477050 219218 477286 219454
rect 477050 218898 477286 219134
rect 473546 186618 474102 187174
rect 480986 194058 481542 194614
rect 477050 183218 477286 183454
rect 477050 182898 477286 183134
rect 473546 150618 474102 151174
rect 480986 158058 481542 158614
rect 477050 147218 477286 147454
rect 477050 146898 477286 147134
rect 473546 114618 474102 115174
rect 480986 122058 481542 122614
rect 477050 111218 477286 111454
rect 477050 110898 477286 111134
rect 473546 78618 474102 79174
rect 480986 86058 481542 86614
rect 477050 75218 477286 75454
rect 477050 74898 477286 75134
rect 473546 42618 474102 43174
rect 480986 50058 481542 50614
rect 477050 39218 477286 39454
rect 477050 38898 477286 39134
rect 473546 6618 474102 7174
rect 473546 -1862 474102 -1306
rect 480986 14058 481542 14614
rect 480986 -3782 481542 -3226
rect 484706 708122 485262 708678
rect 484706 665778 485262 666334
rect 484706 629778 485262 630334
rect 484706 593778 485262 594334
rect 484706 557778 485262 558334
rect 484706 521778 485262 522334
rect 484706 485778 485262 486334
rect 484706 449778 485262 450334
rect 484706 413778 485262 414334
rect 484706 377778 485262 378334
rect 484706 341778 485262 342334
rect 484706 305778 485262 306334
rect 484706 269778 485262 270334
rect 484706 233778 485262 234334
rect 484706 197778 485262 198334
rect 484706 161778 485262 162334
rect 484706 125778 485262 126334
rect 484706 89778 485262 90334
rect 484706 53778 485262 54334
rect 484706 17778 485262 18334
rect 484706 -4742 485262 -4186
rect 488426 709082 488982 709638
rect 488426 669498 488982 670054
rect 488426 633498 488982 634054
rect 488426 597498 488982 598054
rect 488426 561498 488982 562054
rect 488426 525498 488982 526054
rect 488426 489498 488982 490054
rect 488426 453498 488982 454054
rect 488426 417498 488982 418054
rect 488426 381498 488982 382054
rect 492146 710042 492702 710598
rect 492146 673218 492702 673774
rect 492146 637218 492702 637774
rect 492146 601218 492702 601774
rect 492146 565218 492702 565774
rect 492146 529218 492702 529774
rect 492146 493218 492702 493774
rect 492146 457218 492702 457774
rect 492146 421218 492702 421774
rect 492146 385218 492702 385774
rect 495866 711002 496422 711558
rect 495866 676938 496422 677494
rect 495866 640938 496422 641494
rect 495866 604938 496422 605494
rect 495866 568938 496422 569494
rect 495866 532938 496422 533494
rect 495866 496938 496422 497494
rect 495866 460938 496422 461494
rect 495866 424938 496422 425494
rect 495866 388938 496422 389494
rect 488426 345498 488982 346054
rect 495866 352938 496422 353494
rect 492410 330938 492646 331174
rect 492410 330618 492646 330854
rect 488426 309498 488982 310054
rect 495866 316938 496422 317494
rect 492410 294938 492646 295174
rect 492410 294618 492646 294854
rect 488426 273498 488982 274054
rect 495866 280938 496422 281494
rect 492410 258938 492646 259174
rect 492410 258618 492646 258854
rect 488426 237498 488982 238054
rect 495866 244938 496422 245494
rect 492410 222938 492646 223174
rect 492410 222618 492646 222854
rect 488426 201498 488982 202054
rect 495866 208938 496422 209494
rect 492410 186938 492646 187174
rect 492410 186618 492646 186854
rect 488426 165498 488982 166054
rect 495866 172938 496422 173494
rect 492410 150938 492646 151174
rect 492410 150618 492646 150854
rect 488426 129498 488982 130054
rect 495866 136938 496422 137494
rect 492410 114938 492646 115174
rect 492410 114618 492646 114854
rect 488426 93498 488982 94054
rect 495866 100938 496422 101494
rect 492410 78938 492646 79174
rect 492410 78618 492646 78854
rect 488426 57498 488982 58054
rect 495866 64938 496422 65494
rect 492410 42938 492646 43174
rect 492410 42618 492646 42854
rect 488426 21498 488982 22054
rect 495866 28938 496422 29494
rect 492410 6938 492646 7174
rect 492410 6618 492646 6854
rect 488426 -5702 488982 -5146
rect 505826 704282 506382 704838
rect 505826 686898 506382 687454
rect 505826 650898 506382 651454
rect 505826 614898 506382 615454
rect 505826 578898 506382 579454
rect 505826 542898 506382 543454
rect 505826 506898 506382 507454
rect 505826 470898 506382 471454
rect 505826 434898 506382 435454
rect 505826 398898 506382 399454
rect 505826 362898 506382 363454
rect 509546 705242 510102 705798
rect 509546 690618 510102 691174
rect 509546 654618 510102 655174
rect 509546 618618 510102 619174
rect 509546 582618 510102 583174
rect 509546 546618 510102 547174
rect 509546 510618 510102 511174
rect 509546 474618 510102 475174
rect 509546 438618 510102 439174
rect 509546 402618 510102 403174
rect 509546 366618 510102 367174
rect 509546 330618 510102 331174
rect 505826 326898 506382 327454
rect 507770 327218 508006 327454
rect 507770 326898 508006 327134
rect 509546 294618 510102 295174
rect 505826 290898 506382 291454
rect 507770 291218 508006 291454
rect 507770 290898 508006 291134
rect 509546 258618 510102 259174
rect 505826 254898 506382 255454
rect 507770 255218 508006 255454
rect 507770 254898 508006 255134
rect 509546 222618 510102 223174
rect 505826 218898 506382 219454
rect 507770 219218 508006 219454
rect 507770 218898 508006 219134
rect 509546 186618 510102 187174
rect 505826 182898 506382 183454
rect 507770 183218 508006 183454
rect 507770 182898 508006 183134
rect 509546 150618 510102 151174
rect 505826 146898 506382 147454
rect 507770 147218 508006 147454
rect 507770 146898 508006 147134
rect 509546 114618 510102 115174
rect 505826 110898 506382 111454
rect 507770 111218 508006 111454
rect 507770 110898 508006 111134
rect 509546 78618 510102 79174
rect 505826 74898 506382 75454
rect 507770 75218 508006 75454
rect 507770 74898 508006 75134
rect 509546 42618 510102 43174
rect 505826 38898 506382 39454
rect 507770 39218 508006 39454
rect 507770 38898 508006 39134
rect 505826 2898 506382 3454
rect 495866 -7622 496422 -7066
rect 505826 -902 506382 -346
rect 509546 6618 510102 7174
rect 509546 -1862 510102 -1306
rect 513266 706202 513822 706758
rect 513266 694338 513822 694894
rect 513266 658338 513822 658894
rect 513266 622338 513822 622894
rect 513266 586338 513822 586894
rect 513266 550338 513822 550894
rect 513266 514338 513822 514894
rect 513266 478338 513822 478894
rect 513266 442338 513822 442894
rect 513266 406338 513822 406894
rect 513266 370338 513822 370894
rect 513266 334338 513822 334894
rect 513266 298338 513822 298894
rect 513266 262338 513822 262894
rect 513266 226338 513822 226894
rect 513266 190338 513822 190894
rect 513266 154338 513822 154894
rect 513266 118338 513822 118894
rect 513266 82338 513822 82894
rect 513266 46338 513822 46894
rect 513266 10338 513822 10894
rect 516986 707162 517542 707718
rect 516986 698058 517542 698614
rect 516986 662058 517542 662614
rect 516986 626058 517542 626614
rect 516986 590058 517542 590614
rect 516986 554058 517542 554614
rect 516986 518058 517542 518614
rect 516986 482058 517542 482614
rect 516986 446058 517542 446614
rect 516986 410058 517542 410614
rect 516986 374058 517542 374614
rect 516986 338058 517542 338614
rect 516986 302058 517542 302614
rect 516986 266058 517542 266614
rect 516986 230058 517542 230614
rect 516986 194058 517542 194614
rect 516986 158058 517542 158614
rect 516986 122058 517542 122614
rect 516986 86058 517542 86614
rect 516986 50058 517542 50614
rect 516986 14058 517542 14614
rect 513266 -2822 513822 -2266
rect 520706 708122 521262 708678
rect 520706 665778 521262 666334
rect 520706 629778 521262 630334
rect 520706 593778 521262 594334
rect 520706 557778 521262 558334
rect 520706 521778 521262 522334
rect 520706 485778 521262 486334
rect 520706 449778 521262 450334
rect 520706 413778 521262 414334
rect 520706 377778 521262 378334
rect 520706 341778 521262 342334
rect 524426 709082 524982 709638
rect 524426 669498 524982 670054
rect 524426 633498 524982 634054
rect 524426 597498 524982 598054
rect 524426 561498 524982 562054
rect 524426 525498 524982 526054
rect 524426 489498 524982 490054
rect 524426 453498 524982 454054
rect 524426 417498 524982 418054
rect 524426 381498 524982 382054
rect 524426 345498 524982 346054
rect 523130 330938 523366 331174
rect 523130 330618 523366 330854
rect 520706 305778 521262 306334
rect 524426 309498 524982 310054
rect 523130 294938 523366 295174
rect 523130 294618 523366 294854
rect 520706 269778 521262 270334
rect 524426 273498 524982 274054
rect 523130 258938 523366 259174
rect 523130 258618 523366 258854
rect 520706 233778 521262 234334
rect 524426 237498 524982 238054
rect 523130 222938 523366 223174
rect 523130 222618 523366 222854
rect 520706 197778 521262 198334
rect 524426 201498 524982 202054
rect 523130 186938 523366 187174
rect 523130 186618 523366 186854
rect 520706 161778 521262 162334
rect 524426 165498 524982 166054
rect 523130 150938 523366 151174
rect 523130 150618 523366 150854
rect 520706 125778 521262 126334
rect 524426 129498 524982 130054
rect 523130 114938 523366 115174
rect 523130 114618 523366 114854
rect 520706 89778 521262 90334
rect 524426 93498 524982 94054
rect 523130 78938 523366 79174
rect 523130 78618 523366 78854
rect 520706 53778 521262 54334
rect 524426 57498 524982 58054
rect 523130 42938 523366 43174
rect 523130 42618 523366 42854
rect 520706 17778 521262 18334
rect 516986 -3782 517542 -3226
rect 524426 21498 524982 22054
rect 523130 6938 523366 7174
rect 523130 6618 523366 6854
rect 520706 -4742 521262 -4186
rect 528146 710042 528702 710598
rect 528146 673218 528702 673774
rect 528146 637218 528702 637774
rect 528146 601218 528702 601774
rect 528146 565218 528702 565774
rect 528146 529218 528702 529774
rect 528146 493218 528702 493774
rect 528146 457218 528702 457774
rect 528146 421218 528702 421774
rect 528146 385218 528702 385774
rect 528146 349218 528702 349774
rect 528146 313218 528702 313774
rect 528146 277218 528702 277774
rect 528146 241218 528702 241774
rect 528146 205218 528702 205774
rect 528146 169218 528702 169774
rect 528146 133218 528702 133774
rect 528146 97218 528702 97774
rect 528146 61218 528702 61774
rect 528146 25218 528702 25774
rect 524426 -5702 524982 -5146
rect 531866 711002 532422 711558
rect 531866 676938 532422 677494
rect 531866 640938 532422 641494
rect 531866 604938 532422 605494
rect 531866 568938 532422 569494
rect 531866 532938 532422 533494
rect 531866 496938 532422 497494
rect 531866 460938 532422 461494
rect 531866 424938 532422 425494
rect 531866 388938 532422 389494
rect 531866 352938 532422 353494
rect 541826 704282 542382 704838
rect 541826 686898 542382 687454
rect 541826 650898 542382 651454
rect 541826 614898 542382 615454
rect 541826 578898 542382 579454
rect 541826 542898 542382 543454
rect 541826 506898 542382 507454
rect 541826 470898 542382 471454
rect 541826 434898 542382 435454
rect 541826 398898 542382 399454
rect 541826 362898 542382 363454
rect 538490 327218 538726 327454
rect 538490 326898 538726 327134
rect 541826 326898 542382 327454
rect 531866 316938 532422 317494
rect 538490 291218 538726 291454
rect 538490 290898 538726 291134
rect 541826 290898 542382 291454
rect 531866 280938 532422 281494
rect 538490 255218 538726 255454
rect 538490 254898 538726 255134
rect 541826 254898 542382 255454
rect 531866 244938 532422 245494
rect 538490 219218 538726 219454
rect 538490 218898 538726 219134
rect 541826 218898 542382 219454
rect 531866 208938 532422 209494
rect 538490 183218 538726 183454
rect 538490 182898 538726 183134
rect 541826 182898 542382 183454
rect 531866 172938 532422 173494
rect 538490 147218 538726 147454
rect 538490 146898 538726 147134
rect 541826 146898 542382 147454
rect 531866 136938 532422 137494
rect 538490 111218 538726 111454
rect 538490 110898 538726 111134
rect 541826 110898 542382 111454
rect 531866 100938 532422 101494
rect 538490 75218 538726 75454
rect 538490 74898 538726 75134
rect 541826 74898 542382 75454
rect 531866 64938 532422 65494
rect 538490 39218 538726 39454
rect 538490 38898 538726 39134
rect 541826 38898 542382 39454
rect 531866 28938 532422 29494
rect 528146 -6662 528702 -6106
rect 545546 705242 546102 705798
rect 545546 690618 546102 691174
rect 545546 654618 546102 655174
rect 545546 618618 546102 619174
rect 545546 582618 546102 583174
rect 545546 546618 546102 547174
rect 545546 510618 546102 511174
rect 545546 474618 546102 475174
rect 545546 438618 546102 439174
rect 545546 402618 546102 403174
rect 545546 366618 546102 367174
rect 545546 330618 546102 331174
rect 545546 294618 546102 295174
rect 545546 258618 546102 259174
rect 545546 222618 546102 223174
rect 545546 186618 546102 187174
rect 545546 150618 546102 151174
rect 545546 114618 546102 115174
rect 545546 78618 546102 79174
rect 545546 42618 546102 43174
rect 545546 6618 546102 7174
rect 541826 2898 542382 3454
rect 531866 -7622 532422 -7066
rect 541826 -902 542382 -346
rect 549266 706202 549822 706758
rect 549266 694338 549822 694894
rect 549266 658338 549822 658894
rect 549266 622338 549822 622894
rect 549266 586338 549822 586894
rect 549266 550338 549822 550894
rect 549266 514338 549822 514894
rect 549266 478338 549822 478894
rect 549266 442338 549822 442894
rect 549266 406338 549822 406894
rect 549266 370338 549822 370894
rect 549266 334338 549822 334894
rect 549266 298338 549822 298894
rect 549266 262338 549822 262894
rect 549266 226338 549822 226894
rect 549266 190338 549822 190894
rect 549266 154338 549822 154894
rect 549266 118338 549822 118894
rect 549266 82338 549822 82894
rect 549266 46338 549822 46894
rect 549266 10338 549822 10894
rect 545546 -1862 546102 -1306
rect 552986 707162 553542 707718
rect 552986 698058 553542 698614
rect 552986 662058 553542 662614
rect 552986 626058 553542 626614
rect 552986 590058 553542 590614
rect 552986 554058 553542 554614
rect 552986 518058 553542 518614
rect 552986 482058 553542 482614
rect 552986 446058 553542 446614
rect 552986 410058 553542 410614
rect 552986 374058 553542 374614
rect 552986 338058 553542 338614
rect 556706 708122 557262 708678
rect 556706 665778 557262 666334
rect 556706 629778 557262 630334
rect 556706 593778 557262 594334
rect 556706 557778 557262 558334
rect 556706 521778 557262 522334
rect 556706 485778 557262 486334
rect 556706 449778 557262 450334
rect 556706 413778 557262 414334
rect 556706 377778 557262 378334
rect 556706 341778 557262 342334
rect 553850 330938 554086 331174
rect 553850 330618 554086 330854
rect 552986 302058 553542 302614
rect 556706 305778 557262 306334
rect 553850 294938 554086 295174
rect 553850 294618 554086 294854
rect 552986 266058 553542 266614
rect 556706 269778 557262 270334
rect 553850 258938 554086 259174
rect 553850 258618 554086 258854
rect 552986 230058 553542 230614
rect 556706 233778 557262 234334
rect 553850 222938 554086 223174
rect 553850 222618 554086 222854
rect 552986 194058 553542 194614
rect 556706 197778 557262 198334
rect 553850 186938 554086 187174
rect 553850 186618 554086 186854
rect 552986 158058 553542 158614
rect 556706 161778 557262 162334
rect 553850 150938 554086 151174
rect 553850 150618 554086 150854
rect 552986 122058 553542 122614
rect 556706 125778 557262 126334
rect 553850 114938 554086 115174
rect 553850 114618 554086 114854
rect 552986 86058 553542 86614
rect 556706 89778 557262 90334
rect 553850 78938 554086 79174
rect 553850 78618 554086 78854
rect 552986 50058 553542 50614
rect 556706 53778 557262 54334
rect 553850 42938 554086 43174
rect 553850 42618 554086 42854
rect 552986 14058 553542 14614
rect 549266 -2822 549822 -2266
rect 556706 17778 557262 18334
rect 553850 6938 554086 7174
rect 553850 6618 554086 6854
rect 552986 -3782 553542 -3226
rect 560426 709082 560982 709638
rect 560426 669498 560982 670054
rect 560426 633498 560982 634054
rect 560426 597498 560982 598054
rect 560426 561498 560982 562054
rect 560426 525498 560982 526054
rect 560426 489498 560982 490054
rect 560426 453498 560982 454054
rect 560426 417498 560982 418054
rect 560426 381498 560982 382054
rect 560426 345498 560982 346054
rect 560426 309498 560982 310054
rect 560426 273498 560982 274054
rect 560426 237498 560982 238054
rect 560426 201498 560982 202054
rect 560426 165498 560982 166054
rect 560426 129498 560982 130054
rect 560426 93498 560982 94054
rect 560426 57498 560982 58054
rect 560426 21498 560982 22054
rect 556706 -4742 557262 -4186
rect 560426 -5702 560982 -5146
rect 564146 710042 564702 710598
rect 564146 673218 564702 673774
rect 564146 637218 564702 637774
rect 564146 601218 564702 601774
rect 564146 565218 564702 565774
rect 564146 529218 564702 529774
rect 564146 493218 564702 493774
rect 564146 457218 564702 457774
rect 564146 421218 564702 421774
rect 564146 385218 564702 385774
rect 564146 349218 564702 349774
rect 564146 313218 564702 313774
rect 564146 277218 564702 277774
rect 564146 241218 564702 241774
rect 564146 205218 564702 205774
rect 564146 169218 564702 169774
rect 564146 133218 564702 133774
rect 564146 97218 564702 97774
rect 564146 61218 564702 61774
rect 564146 25218 564702 25774
rect 564146 -6662 564702 -6106
rect 567866 711002 568422 711558
rect 567866 676938 568422 677494
rect 567866 640938 568422 641494
rect 567866 604938 568422 605494
rect 567866 568938 568422 569494
rect 567866 532938 568422 533494
rect 567866 496938 568422 497494
rect 567866 460938 568422 461494
rect 567866 424938 568422 425494
rect 567866 388938 568422 389494
rect 567866 352938 568422 353494
rect 577826 704282 578382 704838
rect 577826 686898 578382 687454
rect 577826 650898 578382 651454
rect 577826 614898 578382 615454
rect 577826 578898 578382 579454
rect 577826 542898 578382 543454
rect 577826 506898 578382 507454
rect 577826 470898 578382 471454
rect 577826 434898 578382 435454
rect 577826 398898 578382 399454
rect 577826 362898 578382 363454
rect 569210 327218 569446 327454
rect 569210 326898 569446 327134
rect 567866 316938 568422 317494
rect 577826 326898 578382 327454
rect 569210 291218 569446 291454
rect 569210 290898 569446 291134
rect 567866 280938 568422 281494
rect 577826 290898 578382 291454
rect 569210 255218 569446 255454
rect 569210 254898 569446 255134
rect 567866 244938 568422 245494
rect 577826 254898 578382 255454
rect 569210 219218 569446 219454
rect 569210 218898 569446 219134
rect 567866 208938 568422 209494
rect 577826 218898 578382 219454
rect 569210 183218 569446 183454
rect 569210 182898 569446 183134
rect 567866 172938 568422 173494
rect 577826 182898 578382 183454
rect 569210 147218 569446 147454
rect 569210 146898 569446 147134
rect 567866 136938 568422 137494
rect 577826 146898 578382 147454
rect 569210 111218 569446 111454
rect 569210 110898 569446 111134
rect 567866 100938 568422 101494
rect 577826 110898 578382 111454
rect 569210 75218 569446 75454
rect 569210 74898 569446 75134
rect 577826 74898 578382 75454
rect 567866 64938 568422 65494
rect 569210 39218 569446 39454
rect 569210 38898 569446 39134
rect 577826 38898 578382 39454
rect 567866 28938 568422 29494
rect 567866 -7622 568422 -7066
rect 577826 2898 578382 3454
rect 577826 -902 578382 -346
rect 592062 711002 592618 711558
rect 591102 710042 591658 710598
rect 590142 709082 590698 709638
rect 589182 708122 589738 708678
rect 588222 707162 588778 707718
rect 587262 706202 587818 706758
rect 581546 705242 582102 705798
rect 586302 705242 586858 705798
rect 581546 690618 582102 691174
rect 581546 654618 582102 655174
rect 581546 618618 582102 619174
rect 581546 582618 582102 583174
rect 581546 546618 582102 547174
rect 581546 510618 582102 511174
rect 581546 474618 582102 475174
rect 581546 438618 582102 439174
rect 581546 402618 582102 403174
rect 581546 366618 582102 367174
rect 581546 330618 582102 331174
rect 581546 294618 582102 295174
rect 581546 258618 582102 259174
rect 581546 222618 582102 223174
rect 581546 186618 582102 187174
rect 581546 150618 582102 151174
rect 581546 114618 582102 115174
rect 581546 78618 582102 79174
rect 581546 42618 582102 43174
rect 581546 6618 582102 7174
rect 585342 704282 585898 704838
rect 585342 686898 585898 687454
rect 585342 650898 585898 651454
rect 585342 614898 585898 615454
rect 585342 578898 585898 579454
rect 585342 542898 585898 543454
rect 585342 506898 585898 507454
rect 585342 470898 585898 471454
rect 585342 434898 585898 435454
rect 585342 398898 585898 399454
rect 585342 362898 585898 363454
rect 585342 326898 585898 327454
rect 585342 290898 585898 291454
rect 585342 254898 585898 255454
rect 585342 218898 585898 219454
rect 585342 182898 585898 183454
rect 585342 146898 585898 147454
rect 585342 110898 585898 111454
rect 585342 74898 585898 75454
rect 585342 38898 585898 39454
rect 585342 2898 585898 3454
rect 585342 -902 585898 -346
rect 586302 690618 586858 691174
rect 586302 654618 586858 655174
rect 586302 618618 586858 619174
rect 586302 582618 586858 583174
rect 586302 546618 586858 547174
rect 586302 510618 586858 511174
rect 586302 474618 586858 475174
rect 586302 438618 586858 439174
rect 586302 402618 586858 403174
rect 586302 366618 586858 367174
rect 586302 330618 586858 331174
rect 586302 294618 586858 295174
rect 586302 258618 586858 259174
rect 586302 222618 586858 223174
rect 586302 186618 586858 187174
rect 586302 150618 586858 151174
rect 586302 114618 586858 115174
rect 586302 78618 586858 79174
rect 586302 42618 586858 43174
rect 586302 6618 586858 7174
rect 581546 -1862 582102 -1306
rect 586302 -1862 586858 -1306
rect 587262 694338 587818 694894
rect 587262 658338 587818 658894
rect 587262 622338 587818 622894
rect 587262 586338 587818 586894
rect 587262 550338 587818 550894
rect 587262 514338 587818 514894
rect 587262 478338 587818 478894
rect 587262 442338 587818 442894
rect 587262 406338 587818 406894
rect 587262 370338 587818 370894
rect 587262 334338 587818 334894
rect 587262 298338 587818 298894
rect 587262 262338 587818 262894
rect 587262 226338 587818 226894
rect 587262 190338 587818 190894
rect 587262 154338 587818 154894
rect 587262 118338 587818 118894
rect 587262 82338 587818 82894
rect 587262 46338 587818 46894
rect 587262 10338 587818 10894
rect 587262 -2822 587818 -2266
rect 588222 698058 588778 698614
rect 588222 662058 588778 662614
rect 588222 626058 588778 626614
rect 588222 590058 588778 590614
rect 588222 554058 588778 554614
rect 588222 518058 588778 518614
rect 588222 482058 588778 482614
rect 588222 446058 588778 446614
rect 588222 410058 588778 410614
rect 588222 374058 588778 374614
rect 588222 338058 588778 338614
rect 588222 302058 588778 302614
rect 588222 266058 588778 266614
rect 588222 230058 588778 230614
rect 588222 194058 588778 194614
rect 588222 158058 588778 158614
rect 588222 122058 588778 122614
rect 588222 86058 588778 86614
rect 588222 50058 588778 50614
rect 588222 14058 588778 14614
rect 588222 -3782 588778 -3226
rect 589182 665778 589738 666334
rect 589182 629778 589738 630334
rect 589182 593778 589738 594334
rect 589182 557778 589738 558334
rect 589182 521778 589738 522334
rect 589182 485778 589738 486334
rect 589182 449778 589738 450334
rect 589182 413778 589738 414334
rect 589182 377778 589738 378334
rect 589182 341778 589738 342334
rect 589182 305778 589738 306334
rect 589182 269778 589738 270334
rect 589182 233778 589738 234334
rect 589182 197778 589738 198334
rect 589182 161778 589738 162334
rect 589182 125778 589738 126334
rect 589182 89778 589738 90334
rect 589182 53778 589738 54334
rect 589182 17778 589738 18334
rect 589182 -4742 589738 -4186
rect 590142 669498 590698 670054
rect 590142 633498 590698 634054
rect 590142 597498 590698 598054
rect 590142 561498 590698 562054
rect 590142 525498 590698 526054
rect 590142 489498 590698 490054
rect 590142 453498 590698 454054
rect 590142 417498 590698 418054
rect 590142 381498 590698 382054
rect 590142 345498 590698 346054
rect 590142 309498 590698 310054
rect 590142 273498 590698 274054
rect 590142 237498 590698 238054
rect 590142 201498 590698 202054
rect 590142 165498 590698 166054
rect 590142 129498 590698 130054
rect 590142 93498 590698 94054
rect 590142 57498 590698 58054
rect 590142 21498 590698 22054
rect 590142 -5702 590698 -5146
rect 591102 673218 591658 673774
rect 591102 637218 591658 637774
rect 591102 601218 591658 601774
rect 591102 565218 591658 565774
rect 591102 529218 591658 529774
rect 591102 493218 591658 493774
rect 591102 457218 591658 457774
rect 591102 421218 591658 421774
rect 591102 385218 591658 385774
rect 591102 349218 591658 349774
rect 591102 313218 591658 313774
rect 591102 277218 591658 277774
rect 591102 241218 591658 241774
rect 591102 205218 591658 205774
rect 591102 169218 591658 169774
rect 591102 133218 591658 133774
rect 591102 97218 591658 97774
rect 591102 61218 591658 61774
rect 591102 25218 591658 25774
rect 591102 -6662 591658 -6106
rect 592062 676938 592618 677494
rect 592062 640938 592618 641494
rect 592062 604938 592618 605494
rect 592062 568938 592618 569494
rect 592062 532938 592618 533494
rect 592062 496938 592618 497494
rect 592062 460938 592618 461494
rect 592062 424938 592618 425494
rect 592062 388938 592618 389494
rect 592062 352938 592618 353494
rect 592062 316938 592618 317494
rect 592062 280938 592618 281494
rect 592062 244938 592618 245494
rect 592062 208938 592618 209494
rect 592062 172938 592618 173494
rect 592062 136938 592618 137494
rect 592062 100938 592618 101494
rect 592062 64938 592618 65494
rect 592062 28938 592618 29494
rect 592062 -7622 592618 -7066
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711002 -8694 711558
rect -8138 711002 27866 711558
rect 28422 711002 63866 711558
rect 64422 711002 99866 711558
rect 100422 711002 135866 711558
rect 136422 711002 171866 711558
rect 172422 711002 207866 711558
rect 208422 711002 243866 711558
rect 244422 711002 279866 711558
rect 280422 711002 315866 711558
rect 316422 711002 351866 711558
rect 352422 711002 387866 711558
rect 388422 711002 423866 711558
rect 424422 711002 459866 711558
rect 460422 711002 495866 711558
rect 496422 711002 531866 711558
rect 532422 711002 567866 711558
rect 568422 711002 592062 711558
rect 592618 711002 592650 711558
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710042 -7734 710598
rect -7178 710042 24146 710598
rect 24702 710042 60146 710598
rect 60702 710042 96146 710598
rect 96702 710042 132146 710598
rect 132702 710042 168146 710598
rect 168702 710042 204146 710598
rect 204702 710042 240146 710598
rect 240702 710042 276146 710598
rect 276702 710042 312146 710598
rect 312702 710042 348146 710598
rect 348702 710042 384146 710598
rect 384702 710042 420146 710598
rect 420702 710042 456146 710598
rect 456702 710042 492146 710598
rect 492702 710042 528146 710598
rect 528702 710042 564146 710598
rect 564702 710042 591102 710598
rect 591658 710042 591690 710598
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709082 -6774 709638
rect -6218 709082 20426 709638
rect 20982 709082 56426 709638
rect 56982 709082 92426 709638
rect 92982 709082 128426 709638
rect 128982 709082 164426 709638
rect 164982 709082 200426 709638
rect 200982 709082 236426 709638
rect 236982 709082 272426 709638
rect 272982 709082 308426 709638
rect 308982 709082 344426 709638
rect 344982 709082 380426 709638
rect 380982 709082 416426 709638
rect 416982 709082 452426 709638
rect 452982 709082 488426 709638
rect 488982 709082 524426 709638
rect 524982 709082 560426 709638
rect 560982 709082 590142 709638
rect 590698 709082 590730 709638
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708122 -5814 708678
rect -5258 708122 16706 708678
rect 17262 708122 52706 708678
rect 53262 708122 88706 708678
rect 89262 708122 124706 708678
rect 125262 708122 160706 708678
rect 161262 708122 196706 708678
rect 197262 708122 232706 708678
rect 233262 708122 268706 708678
rect 269262 708122 304706 708678
rect 305262 708122 340706 708678
rect 341262 708122 376706 708678
rect 377262 708122 412706 708678
rect 413262 708122 448706 708678
rect 449262 708122 484706 708678
rect 485262 708122 520706 708678
rect 521262 708122 556706 708678
rect 557262 708122 589182 708678
rect 589738 708122 589770 708678
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707162 -4854 707718
rect -4298 707162 12986 707718
rect 13542 707162 48986 707718
rect 49542 707162 84986 707718
rect 85542 707162 120986 707718
rect 121542 707162 156986 707718
rect 157542 707162 192986 707718
rect 193542 707162 228986 707718
rect 229542 707162 264986 707718
rect 265542 707162 300986 707718
rect 301542 707162 336986 707718
rect 337542 707162 372986 707718
rect 373542 707162 408986 707718
rect 409542 707162 444986 707718
rect 445542 707162 480986 707718
rect 481542 707162 516986 707718
rect 517542 707162 552986 707718
rect 553542 707162 588222 707718
rect 588778 707162 588810 707718
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706202 -3894 706758
rect -3338 706202 9266 706758
rect 9822 706202 45266 706758
rect 45822 706202 81266 706758
rect 81822 706202 117266 706758
rect 117822 706202 153266 706758
rect 153822 706202 189266 706758
rect 189822 706202 225266 706758
rect 225822 706202 261266 706758
rect 261822 706202 297266 706758
rect 297822 706202 333266 706758
rect 333822 706202 369266 706758
rect 369822 706202 405266 706758
rect 405822 706202 441266 706758
rect 441822 706202 477266 706758
rect 477822 706202 513266 706758
rect 513822 706202 549266 706758
rect 549822 706202 587262 706758
rect 587818 706202 587850 706758
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705242 -2934 705798
rect -2378 705242 5546 705798
rect 6102 705242 41546 705798
rect 42102 705242 77546 705798
rect 78102 705242 113546 705798
rect 114102 705242 149546 705798
rect 150102 705242 185546 705798
rect 186102 705242 221546 705798
rect 222102 705242 257546 705798
rect 258102 705242 293546 705798
rect 294102 705242 329546 705798
rect 330102 705242 365546 705798
rect 366102 705242 401546 705798
rect 402102 705242 437546 705798
rect 438102 705242 473546 705798
rect 474102 705242 509546 705798
rect 510102 705242 545546 705798
rect 546102 705242 581546 705798
rect 582102 705242 586302 705798
rect 586858 705242 586890 705798
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704282 -1974 704838
rect -1418 704282 1826 704838
rect 2382 704282 37826 704838
rect 38382 704282 73826 704838
rect 74382 704282 109826 704838
rect 110382 704282 145826 704838
rect 146382 704282 181826 704838
rect 182382 704282 217826 704838
rect 218382 704282 253826 704838
rect 254382 704282 289826 704838
rect 290382 704282 325826 704838
rect 326382 704282 361826 704838
rect 362382 704282 397826 704838
rect 398382 704282 433826 704838
rect 434382 704282 469826 704838
rect 470382 704282 505826 704838
rect 506382 704282 541826 704838
rect 542382 704282 577826 704838
rect 578382 704282 585342 704838
rect 585898 704282 585930 704838
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698058 -4854 698614
rect -4298 698058 12986 698614
rect 13542 698058 48986 698614
rect 49542 698058 84986 698614
rect 85542 698058 120986 698614
rect 121542 698058 156986 698614
rect 157542 698058 192986 698614
rect 193542 698058 228986 698614
rect 229542 698058 264986 698614
rect 265542 698058 300986 698614
rect 301542 698058 336986 698614
rect 337542 698058 372986 698614
rect 373542 698058 408986 698614
rect 409542 698058 444986 698614
rect 445542 698058 480986 698614
rect 481542 698058 516986 698614
rect 517542 698058 552986 698614
rect 553542 698058 588222 698614
rect 588778 698058 592650 698614
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694338 -3894 694894
rect -3338 694338 9266 694894
rect 9822 694338 45266 694894
rect 45822 694338 81266 694894
rect 81822 694338 117266 694894
rect 117822 694338 153266 694894
rect 153822 694338 189266 694894
rect 189822 694338 225266 694894
rect 225822 694338 261266 694894
rect 261822 694338 297266 694894
rect 297822 694338 333266 694894
rect 333822 694338 369266 694894
rect 369822 694338 405266 694894
rect 405822 694338 441266 694894
rect 441822 694338 477266 694894
rect 477822 694338 513266 694894
rect 513822 694338 549266 694894
rect 549822 694338 587262 694894
rect 587818 694338 592650 694894
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690618 -2934 691174
rect -2378 690618 5546 691174
rect 6102 690618 41546 691174
rect 42102 690618 77546 691174
rect 78102 690618 113546 691174
rect 114102 690618 149546 691174
rect 150102 690618 185546 691174
rect 186102 690618 221546 691174
rect 222102 690618 257546 691174
rect 258102 690618 293546 691174
rect 294102 690618 329546 691174
rect 330102 690618 365546 691174
rect 366102 690618 401546 691174
rect 402102 690618 437546 691174
rect 438102 690618 473546 691174
rect 474102 690618 509546 691174
rect 510102 690618 545546 691174
rect 546102 690618 581546 691174
rect 582102 690618 586302 691174
rect 586858 690618 592650 691174
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 686898 -1974 687454
rect -1418 686898 1826 687454
rect 2382 686898 37826 687454
rect 38382 686898 73826 687454
rect 74382 686898 109826 687454
rect 110382 686898 145826 687454
rect 146382 686898 181826 687454
rect 182382 686898 217826 687454
rect 218382 686898 253826 687454
rect 254382 686898 289826 687454
rect 290382 686898 325826 687454
rect 326382 686898 361826 687454
rect 362382 686898 397826 687454
rect 398382 686898 433826 687454
rect 434382 686898 469826 687454
rect 470382 686898 505826 687454
rect 506382 686898 541826 687454
rect 542382 686898 577826 687454
rect 578382 686898 585342 687454
rect 585898 686898 592650 687454
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 676938 -8694 677494
rect -8138 676938 27866 677494
rect 28422 676938 63866 677494
rect 64422 676938 99866 677494
rect 100422 676938 135866 677494
rect 136422 676938 171866 677494
rect 172422 676938 207866 677494
rect 208422 676938 243866 677494
rect 244422 676938 279866 677494
rect 280422 676938 315866 677494
rect 316422 676938 351866 677494
rect 352422 676938 387866 677494
rect 388422 676938 423866 677494
rect 424422 676938 459866 677494
rect 460422 676938 495866 677494
rect 496422 676938 531866 677494
rect 532422 676938 567866 677494
rect 568422 676938 592062 677494
rect 592618 676938 592650 677494
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673218 -7734 673774
rect -7178 673218 24146 673774
rect 24702 673218 60146 673774
rect 60702 673218 96146 673774
rect 96702 673218 132146 673774
rect 132702 673218 168146 673774
rect 168702 673218 204146 673774
rect 204702 673218 240146 673774
rect 240702 673218 276146 673774
rect 276702 673218 312146 673774
rect 312702 673218 348146 673774
rect 348702 673218 384146 673774
rect 384702 673218 420146 673774
rect 420702 673218 456146 673774
rect 456702 673218 492146 673774
rect 492702 673218 528146 673774
rect 528702 673218 564146 673774
rect 564702 673218 591102 673774
rect 591658 673218 592650 673774
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669498 -6774 670054
rect -6218 669498 20426 670054
rect 20982 669498 56426 670054
rect 56982 669498 92426 670054
rect 92982 669498 128426 670054
rect 128982 669498 164426 670054
rect 164982 669498 200426 670054
rect 200982 669498 236426 670054
rect 236982 669498 272426 670054
rect 272982 669498 308426 670054
rect 308982 669498 344426 670054
rect 344982 669498 380426 670054
rect 380982 669498 416426 670054
rect 416982 669498 452426 670054
rect 452982 669498 488426 670054
rect 488982 669498 524426 670054
rect 524982 669498 560426 670054
rect 560982 669498 590142 670054
rect 590698 669498 592650 670054
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 665778 -5814 666334
rect -5258 665778 16706 666334
rect 17262 665778 52706 666334
rect 53262 665778 88706 666334
rect 89262 665778 124706 666334
rect 125262 665778 160706 666334
rect 161262 665778 196706 666334
rect 197262 665778 232706 666334
rect 233262 665778 268706 666334
rect 269262 665778 304706 666334
rect 305262 665778 340706 666334
rect 341262 665778 376706 666334
rect 377262 665778 412706 666334
rect 413262 665778 448706 666334
rect 449262 665778 484706 666334
rect 485262 665778 520706 666334
rect 521262 665778 556706 666334
rect 557262 665778 589182 666334
rect 589738 665778 592650 666334
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662058 -4854 662614
rect -4298 662058 12986 662614
rect 13542 662058 48986 662614
rect 49542 662058 84986 662614
rect 85542 662058 120986 662614
rect 121542 662058 156986 662614
rect 157542 662058 192986 662614
rect 193542 662058 228986 662614
rect 229542 662058 264986 662614
rect 265542 662058 300986 662614
rect 301542 662058 336986 662614
rect 337542 662058 372986 662614
rect 373542 662058 408986 662614
rect 409542 662058 444986 662614
rect 445542 662058 480986 662614
rect 481542 662058 516986 662614
rect 517542 662058 552986 662614
rect 553542 662058 588222 662614
rect 588778 662058 592650 662614
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658338 -3894 658894
rect -3338 658338 9266 658894
rect 9822 658338 45266 658894
rect 45822 658338 81266 658894
rect 81822 658338 117266 658894
rect 117822 658338 153266 658894
rect 153822 658338 189266 658894
rect 189822 658338 225266 658894
rect 225822 658338 261266 658894
rect 261822 658338 297266 658894
rect 297822 658338 333266 658894
rect 333822 658338 369266 658894
rect 369822 658338 405266 658894
rect 405822 658338 441266 658894
rect 441822 658338 477266 658894
rect 477822 658338 513266 658894
rect 513822 658338 549266 658894
rect 549822 658338 587262 658894
rect 587818 658338 592650 658894
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654618 -2934 655174
rect -2378 654618 5546 655174
rect 6102 654618 41546 655174
rect 42102 654618 77546 655174
rect 78102 654618 113546 655174
rect 114102 654618 149546 655174
rect 150102 654618 185546 655174
rect 186102 654618 221546 655174
rect 222102 654618 257546 655174
rect 258102 654618 293546 655174
rect 294102 654618 329546 655174
rect 330102 654618 365546 655174
rect 366102 654618 401546 655174
rect 402102 654618 437546 655174
rect 438102 654618 473546 655174
rect 474102 654618 509546 655174
rect 510102 654618 545546 655174
rect 546102 654618 581546 655174
rect 582102 654618 586302 655174
rect 586858 654618 592650 655174
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 650898 -1974 651454
rect -1418 650898 1826 651454
rect 2382 650898 37826 651454
rect 38382 650898 73826 651454
rect 74382 650898 109826 651454
rect 110382 650898 145826 651454
rect 146382 650898 181826 651454
rect 182382 650898 217826 651454
rect 218382 650898 253826 651454
rect 254382 650898 289826 651454
rect 290382 650898 325826 651454
rect 326382 650898 361826 651454
rect 362382 650898 397826 651454
rect 398382 650898 433826 651454
rect 434382 650898 469826 651454
rect 470382 650898 505826 651454
rect 506382 650898 541826 651454
rect 542382 650898 577826 651454
rect 578382 650898 585342 651454
rect 585898 650898 592650 651454
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 640938 -8694 641494
rect -8138 640938 27866 641494
rect 28422 640938 63866 641494
rect 64422 640938 99866 641494
rect 100422 640938 135866 641494
rect 136422 640938 171866 641494
rect 172422 640938 207866 641494
rect 208422 640938 243866 641494
rect 244422 640938 279866 641494
rect 280422 640938 315866 641494
rect 316422 640938 351866 641494
rect 352422 640938 387866 641494
rect 388422 640938 423866 641494
rect 424422 640938 459866 641494
rect 460422 640938 495866 641494
rect 496422 640938 531866 641494
rect 532422 640938 567866 641494
rect 568422 640938 592062 641494
rect 592618 640938 592650 641494
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637218 -7734 637774
rect -7178 637218 24146 637774
rect 24702 637218 60146 637774
rect 60702 637218 96146 637774
rect 96702 637218 132146 637774
rect 132702 637218 168146 637774
rect 168702 637218 204146 637774
rect 204702 637218 240146 637774
rect 240702 637218 276146 637774
rect 276702 637218 312146 637774
rect 312702 637218 348146 637774
rect 348702 637218 384146 637774
rect 384702 637218 420146 637774
rect 420702 637218 456146 637774
rect 456702 637218 492146 637774
rect 492702 637218 528146 637774
rect 528702 637218 564146 637774
rect 564702 637218 591102 637774
rect 591658 637218 592650 637774
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633498 -6774 634054
rect -6218 633498 20426 634054
rect 20982 633498 56426 634054
rect 56982 633498 92426 634054
rect 92982 633498 128426 634054
rect 128982 633498 164426 634054
rect 164982 633498 200426 634054
rect 200982 633498 236426 634054
rect 236982 633498 272426 634054
rect 272982 633498 308426 634054
rect 308982 633498 344426 634054
rect 344982 633498 380426 634054
rect 380982 633498 416426 634054
rect 416982 633498 452426 634054
rect 452982 633498 488426 634054
rect 488982 633498 524426 634054
rect 524982 633498 560426 634054
rect 560982 633498 590142 634054
rect 590698 633498 592650 634054
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 629778 -5814 630334
rect -5258 629778 16706 630334
rect 17262 629778 52706 630334
rect 53262 629778 88706 630334
rect 89262 629778 124706 630334
rect 125262 629778 160706 630334
rect 161262 629778 196706 630334
rect 197262 629778 232706 630334
rect 233262 629778 268706 630334
rect 269262 629778 304706 630334
rect 305262 629778 340706 630334
rect 341262 629778 376706 630334
rect 377262 629778 412706 630334
rect 413262 629778 448706 630334
rect 449262 629778 484706 630334
rect 485262 629778 520706 630334
rect 521262 629778 556706 630334
rect 557262 629778 589182 630334
rect 589738 629778 592650 630334
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626058 -4854 626614
rect -4298 626058 12986 626614
rect 13542 626058 48986 626614
rect 49542 626058 84986 626614
rect 85542 626058 120986 626614
rect 121542 626058 156986 626614
rect 157542 626058 192986 626614
rect 193542 626058 228986 626614
rect 229542 626058 264986 626614
rect 265542 626058 300986 626614
rect 301542 626058 336986 626614
rect 337542 626058 372986 626614
rect 373542 626058 408986 626614
rect 409542 626058 444986 626614
rect 445542 626058 480986 626614
rect 481542 626058 516986 626614
rect 517542 626058 552986 626614
rect 553542 626058 588222 626614
rect 588778 626058 592650 626614
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622338 -3894 622894
rect -3338 622338 9266 622894
rect 9822 622338 45266 622894
rect 45822 622338 81266 622894
rect 81822 622338 117266 622894
rect 117822 622338 153266 622894
rect 153822 622338 189266 622894
rect 189822 622338 225266 622894
rect 225822 622338 261266 622894
rect 261822 622338 297266 622894
rect 297822 622338 333266 622894
rect 333822 622338 369266 622894
rect 369822 622338 405266 622894
rect 405822 622338 441266 622894
rect 441822 622338 477266 622894
rect 477822 622338 513266 622894
rect 513822 622338 549266 622894
rect 549822 622338 587262 622894
rect 587818 622338 592650 622894
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618618 -2934 619174
rect -2378 618618 5546 619174
rect 6102 618618 41546 619174
rect 42102 618618 77546 619174
rect 78102 618618 113546 619174
rect 114102 618618 149546 619174
rect 150102 618618 185546 619174
rect 186102 618618 221546 619174
rect 222102 618618 257546 619174
rect 258102 618618 293546 619174
rect 294102 618618 329546 619174
rect 330102 618618 365546 619174
rect 366102 618618 401546 619174
rect 402102 618618 437546 619174
rect 438102 618618 473546 619174
rect 474102 618618 509546 619174
rect 510102 618618 545546 619174
rect 546102 618618 581546 619174
rect 582102 618618 586302 619174
rect 586858 618618 592650 619174
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 614898 -1974 615454
rect -1418 614898 1826 615454
rect 2382 614898 37826 615454
rect 38382 614898 73826 615454
rect 74382 614898 109826 615454
rect 110382 614898 145826 615454
rect 146382 614898 181826 615454
rect 182382 614898 217826 615454
rect 218382 614898 253826 615454
rect 254382 614898 289826 615454
rect 290382 614898 325826 615454
rect 326382 614898 361826 615454
rect 362382 614898 397826 615454
rect 398382 614898 433826 615454
rect 434382 614898 469826 615454
rect 470382 614898 505826 615454
rect 506382 614898 541826 615454
rect 542382 614898 577826 615454
rect 578382 614898 585342 615454
rect 585898 614898 592650 615454
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 604938 -8694 605494
rect -8138 604938 27866 605494
rect 28422 604938 63866 605494
rect 64422 604938 99866 605494
rect 100422 604938 135866 605494
rect 136422 604938 171866 605494
rect 172422 604938 207866 605494
rect 208422 604938 243866 605494
rect 244422 604938 279866 605494
rect 280422 604938 315866 605494
rect 316422 604938 351866 605494
rect 352422 604938 387866 605494
rect 388422 604938 423866 605494
rect 424422 604938 459866 605494
rect 460422 604938 495866 605494
rect 496422 604938 531866 605494
rect 532422 604938 567866 605494
rect 568422 604938 592062 605494
rect 592618 604938 592650 605494
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601218 -7734 601774
rect -7178 601218 24146 601774
rect 24702 601218 60146 601774
rect 60702 601218 96146 601774
rect 96702 601218 132146 601774
rect 132702 601218 168146 601774
rect 168702 601218 204146 601774
rect 204702 601218 240146 601774
rect 240702 601218 276146 601774
rect 276702 601218 312146 601774
rect 312702 601218 348146 601774
rect 348702 601218 384146 601774
rect 384702 601218 420146 601774
rect 420702 601218 456146 601774
rect 456702 601218 492146 601774
rect 492702 601218 528146 601774
rect 528702 601218 564146 601774
rect 564702 601218 591102 601774
rect 591658 601218 592650 601774
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597498 -6774 598054
rect -6218 597498 20426 598054
rect 20982 597498 56426 598054
rect 56982 597498 92426 598054
rect 92982 597498 128426 598054
rect 128982 597498 164426 598054
rect 164982 597498 200426 598054
rect 200982 597498 236426 598054
rect 236982 597498 272426 598054
rect 272982 597498 308426 598054
rect 308982 597498 344426 598054
rect 344982 597498 380426 598054
rect 380982 597498 416426 598054
rect 416982 597498 452426 598054
rect 452982 597498 488426 598054
rect 488982 597498 524426 598054
rect 524982 597498 560426 598054
rect 560982 597498 590142 598054
rect 590698 597498 592650 598054
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 593778 -5814 594334
rect -5258 593778 16706 594334
rect 17262 593778 52706 594334
rect 53262 593778 88706 594334
rect 89262 593778 124706 594334
rect 125262 593778 160706 594334
rect 161262 593778 196706 594334
rect 197262 593778 232706 594334
rect 233262 593778 268706 594334
rect 269262 593778 304706 594334
rect 305262 593778 340706 594334
rect 341262 593778 376706 594334
rect 377262 593778 412706 594334
rect 413262 593778 448706 594334
rect 449262 593778 484706 594334
rect 485262 593778 520706 594334
rect 521262 593778 556706 594334
rect 557262 593778 589182 594334
rect 589738 593778 592650 594334
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590058 -4854 590614
rect -4298 590058 12986 590614
rect 13542 590058 48986 590614
rect 49542 590058 84986 590614
rect 85542 590058 120986 590614
rect 121542 590058 156986 590614
rect 157542 590058 192986 590614
rect 193542 590058 228986 590614
rect 229542 590058 264986 590614
rect 265542 590058 300986 590614
rect 301542 590058 336986 590614
rect 337542 590058 372986 590614
rect 373542 590058 408986 590614
rect 409542 590058 444986 590614
rect 445542 590058 480986 590614
rect 481542 590058 516986 590614
rect 517542 590058 552986 590614
rect 553542 590058 588222 590614
rect 588778 590058 592650 590614
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586338 -3894 586894
rect -3338 586338 9266 586894
rect 9822 586338 45266 586894
rect 45822 586338 81266 586894
rect 81822 586338 117266 586894
rect 117822 586338 153266 586894
rect 153822 586338 189266 586894
rect 189822 586338 225266 586894
rect 225822 586338 261266 586894
rect 261822 586338 297266 586894
rect 297822 586338 333266 586894
rect 333822 586338 369266 586894
rect 369822 586338 405266 586894
rect 405822 586338 441266 586894
rect 441822 586338 477266 586894
rect 477822 586338 513266 586894
rect 513822 586338 549266 586894
rect 549822 586338 587262 586894
rect 587818 586338 592650 586894
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582618 -2934 583174
rect -2378 582618 5546 583174
rect 6102 582618 41546 583174
rect 42102 582618 77546 583174
rect 78102 582618 113546 583174
rect 114102 582618 149546 583174
rect 150102 582618 185546 583174
rect 186102 582618 221546 583174
rect 222102 582618 257546 583174
rect 258102 582618 293546 583174
rect 294102 582618 329546 583174
rect 330102 582618 365546 583174
rect 366102 582618 401546 583174
rect 402102 582618 437546 583174
rect 438102 582618 473546 583174
rect 474102 582618 509546 583174
rect 510102 582618 545546 583174
rect 546102 582618 581546 583174
rect 582102 582618 586302 583174
rect 586858 582618 592650 583174
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 578898 -1974 579454
rect -1418 578898 1826 579454
rect 2382 578898 37826 579454
rect 38382 578898 73826 579454
rect 74382 578898 109826 579454
rect 110382 578898 145826 579454
rect 146382 578898 181826 579454
rect 182382 578898 217826 579454
rect 218382 578898 253826 579454
rect 254382 578898 289826 579454
rect 290382 578898 325826 579454
rect 326382 578898 361826 579454
rect 362382 578898 397826 579454
rect 398382 578898 433826 579454
rect 434382 578898 469826 579454
rect 470382 578898 505826 579454
rect 506382 578898 541826 579454
rect 542382 578898 577826 579454
rect 578382 578898 585342 579454
rect 585898 578898 592650 579454
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 568938 -8694 569494
rect -8138 568938 27866 569494
rect 28422 568938 63866 569494
rect 64422 568938 99866 569494
rect 100422 568938 135866 569494
rect 136422 568938 171866 569494
rect 172422 568938 207866 569494
rect 208422 568938 243866 569494
rect 244422 568938 279866 569494
rect 280422 568938 315866 569494
rect 316422 568938 351866 569494
rect 352422 568938 387866 569494
rect 388422 568938 423866 569494
rect 424422 568938 459866 569494
rect 460422 568938 495866 569494
rect 496422 568938 531866 569494
rect 532422 568938 567866 569494
rect 568422 568938 592062 569494
rect 592618 568938 592650 569494
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565218 -7734 565774
rect -7178 565218 24146 565774
rect 24702 565218 60146 565774
rect 60702 565218 96146 565774
rect 96702 565218 132146 565774
rect 132702 565218 168146 565774
rect 168702 565218 204146 565774
rect 204702 565218 240146 565774
rect 240702 565218 276146 565774
rect 276702 565218 312146 565774
rect 312702 565218 348146 565774
rect 348702 565218 384146 565774
rect 384702 565218 420146 565774
rect 420702 565218 456146 565774
rect 456702 565218 492146 565774
rect 492702 565218 528146 565774
rect 528702 565218 564146 565774
rect 564702 565218 591102 565774
rect 591658 565218 592650 565774
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561498 -6774 562054
rect -6218 561498 20426 562054
rect 20982 561498 56426 562054
rect 56982 561498 92426 562054
rect 92982 561498 128426 562054
rect 128982 561498 164426 562054
rect 164982 561498 200426 562054
rect 200982 561498 236426 562054
rect 236982 561498 272426 562054
rect 272982 561498 308426 562054
rect 308982 561498 344426 562054
rect 344982 561498 380426 562054
rect 380982 561498 416426 562054
rect 416982 561498 452426 562054
rect 452982 561498 488426 562054
rect 488982 561498 524426 562054
rect 524982 561498 560426 562054
rect 560982 561498 590142 562054
rect 590698 561498 592650 562054
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 557778 -5814 558334
rect -5258 557778 16706 558334
rect 17262 557778 52706 558334
rect 53262 557778 88706 558334
rect 89262 557778 124706 558334
rect 125262 557778 160706 558334
rect 161262 557778 196706 558334
rect 197262 557778 232706 558334
rect 233262 557778 268706 558334
rect 269262 557778 304706 558334
rect 305262 557778 340706 558334
rect 341262 557778 376706 558334
rect 377262 557778 412706 558334
rect 413262 557778 448706 558334
rect 449262 557778 484706 558334
rect 485262 557778 520706 558334
rect 521262 557778 556706 558334
rect 557262 557778 589182 558334
rect 589738 557778 592650 558334
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554058 -4854 554614
rect -4298 554058 12986 554614
rect 13542 554058 48986 554614
rect 49542 554058 84986 554614
rect 85542 554058 120986 554614
rect 121542 554058 156986 554614
rect 157542 554058 192986 554614
rect 193542 554058 228986 554614
rect 229542 554058 264986 554614
rect 265542 554058 300986 554614
rect 301542 554058 336986 554614
rect 337542 554058 372986 554614
rect 373542 554058 408986 554614
rect 409542 554058 444986 554614
rect 445542 554058 480986 554614
rect 481542 554058 516986 554614
rect 517542 554058 552986 554614
rect 553542 554058 588222 554614
rect 588778 554058 592650 554614
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550338 -3894 550894
rect -3338 550338 9266 550894
rect 9822 550338 45266 550894
rect 45822 550338 81266 550894
rect 81822 550338 117266 550894
rect 117822 550338 153266 550894
rect 153822 550338 189266 550894
rect 189822 550338 225266 550894
rect 225822 550338 261266 550894
rect 261822 550338 297266 550894
rect 297822 550338 333266 550894
rect 333822 550338 369266 550894
rect 369822 550338 405266 550894
rect 405822 550338 441266 550894
rect 441822 550338 477266 550894
rect 477822 550338 513266 550894
rect 513822 550338 549266 550894
rect 549822 550338 587262 550894
rect 587818 550338 592650 550894
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546618 -2934 547174
rect -2378 546618 5546 547174
rect 6102 546618 41546 547174
rect 42102 546618 77546 547174
rect 78102 546618 113546 547174
rect 114102 546618 149546 547174
rect 150102 546618 185546 547174
rect 186102 546618 221546 547174
rect 222102 546618 257546 547174
rect 258102 546618 293546 547174
rect 294102 546618 329546 547174
rect 330102 546618 365546 547174
rect 366102 546618 401546 547174
rect 402102 546618 437546 547174
rect 438102 546618 473546 547174
rect 474102 546618 509546 547174
rect 510102 546618 545546 547174
rect 546102 546618 581546 547174
rect 582102 546618 586302 547174
rect 586858 546618 592650 547174
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 542898 -1974 543454
rect -1418 542898 1826 543454
rect 2382 542898 37826 543454
rect 38382 542898 73826 543454
rect 74382 542898 109826 543454
rect 110382 542898 145826 543454
rect 146382 542898 181826 543454
rect 182382 542898 217826 543454
rect 218382 542898 253826 543454
rect 254382 542898 289826 543454
rect 290382 542898 325826 543454
rect 326382 542898 361826 543454
rect 362382 542898 397826 543454
rect 398382 542898 433826 543454
rect 434382 542898 469826 543454
rect 470382 542898 505826 543454
rect 506382 542898 541826 543454
rect 542382 542898 577826 543454
rect 578382 542898 585342 543454
rect 585898 542898 592650 543454
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 532938 -8694 533494
rect -8138 532938 27866 533494
rect 28422 532938 63866 533494
rect 64422 532938 99866 533494
rect 100422 532938 135866 533494
rect 136422 532938 171866 533494
rect 172422 532938 207866 533494
rect 208422 532938 243866 533494
rect 244422 532938 279866 533494
rect 280422 532938 315866 533494
rect 316422 532938 351866 533494
rect 352422 532938 387866 533494
rect 388422 532938 423866 533494
rect 424422 532938 459866 533494
rect 460422 532938 495866 533494
rect 496422 532938 531866 533494
rect 532422 532938 567866 533494
rect 568422 532938 592062 533494
rect 592618 532938 592650 533494
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529218 -7734 529774
rect -7178 529218 24146 529774
rect 24702 529218 60146 529774
rect 60702 529218 96146 529774
rect 96702 529218 132146 529774
rect 132702 529218 168146 529774
rect 168702 529218 204146 529774
rect 204702 529218 240146 529774
rect 240702 529218 276146 529774
rect 276702 529218 312146 529774
rect 312702 529218 348146 529774
rect 348702 529218 384146 529774
rect 384702 529218 420146 529774
rect 420702 529218 456146 529774
rect 456702 529218 492146 529774
rect 492702 529218 528146 529774
rect 528702 529218 564146 529774
rect 564702 529218 591102 529774
rect 591658 529218 592650 529774
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525498 -6774 526054
rect -6218 525498 20426 526054
rect 20982 525498 56426 526054
rect 56982 525498 92426 526054
rect 92982 525498 128426 526054
rect 128982 525498 164426 526054
rect 164982 525498 200426 526054
rect 200982 525498 236426 526054
rect 236982 525498 272426 526054
rect 272982 525498 308426 526054
rect 308982 525498 344426 526054
rect 344982 525498 380426 526054
rect 380982 525498 416426 526054
rect 416982 525498 452426 526054
rect 452982 525498 488426 526054
rect 488982 525498 524426 526054
rect 524982 525498 560426 526054
rect 560982 525498 590142 526054
rect 590698 525498 592650 526054
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 521778 -5814 522334
rect -5258 521778 16706 522334
rect 17262 521778 52706 522334
rect 53262 521778 88706 522334
rect 89262 521778 124706 522334
rect 125262 521778 160706 522334
rect 161262 521778 196706 522334
rect 197262 521778 232706 522334
rect 233262 521778 268706 522334
rect 269262 521778 304706 522334
rect 305262 521778 340706 522334
rect 341262 521778 376706 522334
rect 377262 521778 412706 522334
rect 413262 521778 448706 522334
rect 449262 521778 484706 522334
rect 485262 521778 520706 522334
rect 521262 521778 556706 522334
rect 557262 521778 589182 522334
rect 589738 521778 592650 522334
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518058 -4854 518614
rect -4298 518058 12986 518614
rect 13542 518058 48986 518614
rect 49542 518058 84986 518614
rect 85542 518058 120986 518614
rect 121542 518058 156986 518614
rect 157542 518058 192986 518614
rect 193542 518058 228986 518614
rect 229542 518058 264986 518614
rect 265542 518058 300986 518614
rect 301542 518058 336986 518614
rect 337542 518058 372986 518614
rect 373542 518058 408986 518614
rect 409542 518058 444986 518614
rect 445542 518058 480986 518614
rect 481542 518058 516986 518614
rect 517542 518058 552986 518614
rect 553542 518058 588222 518614
rect 588778 518058 592650 518614
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514338 -3894 514894
rect -3338 514338 9266 514894
rect 9822 514338 45266 514894
rect 45822 514338 81266 514894
rect 81822 514338 117266 514894
rect 117822 514338 153266 514894
rect 153822 514338 189266 514894
rect 189822 514338 225266 514894
rect 225822 514338 261266 514894
rect 261822 514338 297266 514894
rect 297822 514338 333266 514894
rect 333822 514338 369266 514894
rect 369822 514338 405266 514894
rect 405822 514338 441266 514894
rect 441822 514338 477266 514894
rect 477822 514338 513266 514894
rect 513822 514338 549266 514894
rect 549822 514338 587262 514894
rect 587818 514338 592650 514894
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510618 -2934 511174
rect -2378 510618 5546 511174
rect 6102 510618 41546 511174
rect 42102 510618 77546 511174
rect 78102 510618 113546 511174
rect 114102 510618 149546 511174
rect 150102 510618 185546 511174
rect 186102 510618 221546 511174
rect 222102 510618 257546 511174
rect 258102 510618 293546 511174
rect 294102 510618 329546 511174
rect 330102 510618 365546 511174
rect 366102 510618 401546 511174
rect 402102 510618 437546 511174
rect 438102 510618 473546 511174
rect 474102 510618 509546 511174
rect 510102 510618 545546 511174
rect 546102 510618 581546 511174
rect 582102 510618 586302 511174
rect 586858 510618 592650 511174
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 506898 -1974 507454
rect -1418 506898 1826 507454
rect 2382 506898 37826 507454
rect 38382 506898 73826 507454
rect 74382 506898 109826 507454
rect 110382 506898 145826 507454
rect 146382 506898 181826 507454
rect 182382 506898 217826 507454
rect 218382 506898 253826 507454
rect 254382 506898 289826 507454
rect 290382 506898 325826 507454
rect 326382 506898 361826 507454
rect 362382 506898 397826 507454
rect 398382 506898 433826 507454
rect 434382 506898 469826 507454
rect 470382 506898 505826 507454
rect 506382 506898 541826 507454
rect 542382 506898 577826 507454
rect 578382 506898 585342 507454
rect 585898 506898 592650 507454
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 496938 -8694 497494
rect -8138 496938 27866 497494
rect 28422 496938 63866 497494
rect 64422 496938 99866 497494
rect 100422 496938 135866 497494
rect 136422 496938 171866 497494
rect 172422 496938 207866 497494
rect 208422 496938 243866 497494
rect 244422 496938 279866 497494
rect 280422 496938 315866 497494
rect 316422 496938 351866 497494
rect 352422 496938 387866 497494
rect 388422 496938 423866 497494
rect 424422 496938 459866 497494
rect 460422 496938 495866 497494
rect 496422 496938 531866 497494
rect 532422 496938 567866 497494
rect 568422 496938 592062 497494
rect 592618 496938 592650 497494
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493218 -7734 493774
rect -7178 493218 24146 493774
rect 24702 493218 60146 493774
rect 60702 493218 96146 493774
rect 96702 493218 132146 493774
rect 132702 493218 168146 493774
rect 168702 493218 204146 493774
rect 204702 493218 240146 493774
rect 240702 493218 276146 493774
rect 276702 493218 312146 493774
rect 312702 493218 348146 493774
rect 348702 493218 384146 493774
rect 384702 493218 420146 493774
rect 420702 493218 456146 493774
rect 456702 493218 492146 493774
rect 492702 493218 528146 493774
rect 528702 493218 564146 493774
rect 564702 493218 591102 493774
rect 591658 493218 592650 493774
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489498 -6774 490054
rect -6218 489498 20426 490054
rect 20982 489498 56426 490054
rect 56982 489498 92426 490054
rect 92982 489498 128426 490054
rect 128982 489498 164426 490054
rect 164982 489498 200426 490054
rect 200982 489498 236426 490054
rect 236982 489498 272426 490054
rect 272982 489498 308426 490054
rect 308982 489498 344426 490054
rect 344982 489498 380426 490054
rect 380982 489498 416426 490054
rect 416982 489498 452426 490054
rect 452982 489498 488426 490054
rect 488982 489498 524426 490054
rect 524982 489498 560426 490054
rect 560982 489498 590142 490054
rect 590698 489498 592650 490054
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 485778 -5814 486334
rect -5258 485778 16706 486334
rect 17262 485778 52706 486334
rect 53262 485778 88706 486334
rect 89262 485778 124706 486334
rect 125262 485778 160706 486334
rect 161262 485778 196706 486334
rect 197262 485778 232706 486334
rect 233262 485778 268706 486334
rect 269262 485778 304706 486334
rect 305262 485778 340706 486334
rect 341262 485778 376706 486334
rect 377262 485778 412706 486334
rect 413262 485778 448706 486334
rect 449262 485778 484706 486334
rect 485262 485778 520706 486334
rect 521262 485778 556706 486334
rect 557262 485778 589182 486334
rect 589738 485778 592650 486334
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482058 -4854 482614
rect -4298 482058 12986 482614
rect 13542 482058 48986 482614
rect 49542 482058 84986 482614
rect 85542 482058 120986 482614
rect 121542 482058 156986 482614
rect 157542 482058 192986 482614
rect 193542 482058 228986 482614
rect 229542 482058 264986 482614
rect 265542 482058 300986 482614
rect 301542 482058 336986 482614
rect 337542 482058 372986 482614
rect 373542 482058 408986 482614
rect 409542 482058 444986 482614
rect 445542 482058 480986 482614
rect 481542 482058 516986 482614
rect 517542 482058 552986 482614
rect 553542 482058 588222 482614
rect 588778 482058 592650 482614
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478338 -3894 478894
rect -3338 478338 9266 478894
rect 9822 478338 45266 478894
rect 45822 478338 81266 478894
rect 81822 478338 117266 478894
rect 117822 478338 153266 478894
rect 153822 478338 189266 478894
rect 189822 478338 225266 478894
rect 225822 478338 261266 478894
rect 261822 478338 297266 478894
rect 297822 478338 333266 478894
rect 333822 478338 369266 478894
rect 369822 478338 405266 478894
rect 405822 478338 441266 478894
rect 441822 478338 477266 478894
rect 477822 478338 513266 478894
rect 513822 478338 549266 478894
rect 549822 478338 587262 478894
rect 587818 478338 592650 478894
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474618 -2934 475174
rect -2378 474618 5546 475174
rect 6102 474618 41546 475174
rect 42102 474618 77546 475174
rect 78102 474618 113546 475174
rect 114102 474618 149546 475174
rect 150102 474618 185546 475174
rect 186102 474618 221546 475174
rect 222102 474618 257546 475174
rect 258102 474618 293546 475174
rect 294102 474618 329546 475174
rect 330102 474618 365546 475174
rect 366102 474618 401546 475174
rect 402102 474618 437546 475174
rect 438102 474618 473546 475174
rect 474102 474618 509546 475174
rect 510102 474618 545546 475174
rect 546102 474618 581546 475174
rect 582102 474618 586302 475174
rect 586858 474618 592650 475174
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 470898 -1974 471454
rect -1418 470898 1826 471454
rect 2382 470898 37826 471454
rect 38382 470898 73826 471454
rect 74382 470898 109826 471454
rect 110382 470898 145826 471454
rect 146382 470898 181826 471454
rect 182382 470898 217826 471454
rect 218382 470898 253826 471454
rect 254382 470898 289826 471454
rect 290382 470898 325826 471454
rect 326382 470898 361826 471454
rect 362382 470898 397826 471454
rect 398382 470898 433826 471454
rect 434382 470898 469826 471454
rect 470382 470898 505826 471454
rect 506382 470898 541826 471454
rect 542382 470898 577826 471454
rect 578382 470898 585342 471454
rect 585898 470898 592650 471454
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 460938 -8694 461494
rect -8138 460938 27866 461494
rect 28422 460938 63866 461494
rect 64422 460938 99866 461494
rect 100422 460938 135866 461494
rect 136422 460938 171866 461494
rect 172422 460938 207866 461494
rect 208422 460938 243866 461494
rect 244422 460938 279866 461494
rect 280422 460938 315866 461494
rect 316422 460938 351866 461494
rect 352422 460938 387866 461494
rect 388422 460938 423866 461494
rect 424422 460938 459866 461494
rect 460422 460938 495866 461494
rect 496422 460938 531866 461494
rect 532422 460938 567866 461494
rect 568422 460938 592062 461494
rect 592618 460938 592650 461494
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457218 -7734 457774
rect -7178 457218 24146 457774
rect 24702 457218 60146 457774
rect 60702 457218 96146 457774
rect 96702 457218 132146 457774
rect 132702 457218 168146 457774
rect 168702 457218 204146 457774
rect 204702 457218 240146 457774
rect 240702 457218 276146 457774
rect 276702 457218 312146 457774
rect 312702 457218 348146 457774
rect 348702 457218 384146 457774
rect 384702 457218 420146 457774
rect 420702 457218 456146 457774
rect 456702 457218 492146 457774
rect 492702 457218 528146 457774
rect 528702 457218 564146 457774
rect 564702 457218 591102 457774
rect 591658 457218 592650 457774
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453498 -6774 454054
rect -6218 453498 20426 454054
rect 20982 453498 56426 454054
rect 56982 453498 92426 454054
rect 92982 453498 128426 454054
rect 128982 453498 164426 454054
rect 164982 453498 200426 454054
rect 200982 453498 236426 454054
rect 236982 453498 272426 454054
rect 272982 453498 308426 454054
rect 308982 453498 344426 454054
rect 344982 453498 380426 454054
rect 380982 453498 416426 454054
rect 416982 453498 452426 454054
rect 452982 453498 488426 454054
rect 488982 453498 524426 454054
rect 524982 453498 560426 454054
rect 560982 453498 590142 454054
rect 590698 453498 592650 454054
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 449778 -5814 450334
rect -5258 449778 16706 450334
rect 17262 449778 52706 450334
rect 53262 449778 88706 450334
rect 89262 449778 124706 450334
rect 125262 449778 160706 450334
rect 161262 449778 196706 450334
rect 197262 449778 232706 450334
rect 233262 449778 268706 450334
rect 269262 449778 304706 450334
rect 305262 449778 340706 450334
rect 341262 449778 376706 450334
rect 377262 449778 412706 450334
rect 413262 449778 448706 450334
rect 449262 449778 484706 450334
rect 485262 449778 520706 450334
rect 521262 449778 556706 450334
rect 557262 449778 589182 450334
rect 589738 449778 592650 450334
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446058 -4854 446614
rect -4298 446058 12986 446614
rect 13542 446058 48986 446614
rect 49542 446058 84986 446614
rect 85542 446058 120986 446614
rect 121542 446058 156986 446614
rect 157542 446058 192986 446614
rect 193542 446058 228986 446614
rect 229542 446058 264986 446614
rect 265542 446058 300986 446614
rect 301542 446058 336986 446614
rect 337542 446058 372986 446614
rect 373542 446058 408986 446614
rect 409542 446058 444986 446614
rect 445542 446058 480986 446614
rect 481542 446058 516986 446614
rect 517542 446058 552986 446614
rect 553542 446058 588222 446614
rect 588778 446058 592650 446614
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442338 -3894 442894
rect -3338 442338 9266 442894
rect 9822 442338 45266 442894
rect 45822 442338 81266 442894
rect 81822 442338 117266 442894
rect 117822 442338 153266 442894
rect 153822 442338 189266 442894
rect 189822 442338 225266 442894
rect 225822 442338 261266 442894
rect 261822 442338 297266 442894
rect 297822 442338 333266 442894
rect 333822 442338 369266 442894
rect 369822 442338 405266 442894
rect 405822 442338 441266 442894
rect 441822 442338 477266 442894
rect 477822 442338 513266 442894
rect 513822 442338 549266 442894
rect 549822 442338 587262 442894
rect 587818 442338 592650 442894
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438618 -2934 439174
rect -2378 438618 5546 439174
rect 6102 438618 41546 439174
rect 42102 438618 77546 439174
rect 78102 438618 113546 439174
rect 114102 438618 149546 439174
rect 150102 438618 185546 439174
rect 186102 438618 221546 439174
rect 222102 438618 257546 439174
rect 258102 438618 293546 439174
rect 294102 438618 329546 439174
rect 330102 438618 365546 439174
rect 366102 438618 401546 439174
rect 402102 438618 437546 439174
rect 438102 438618 473546 439174
rect 474102 438618 509546 439174
rect 510102 438618 545546 439174
rect 546102 438618 581546 439174
rect 582102 438618 586302 439174
rect 586858 438618 592650 439174
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 434898 -1974 435454
rect -1418 434898 1826 435454
rect 2382 434898 37826 435454
rect 38382 434898 73826 435454
rect 74382 434898 109826 435454
rect 110382 434898 145826 435454
rect 146382 434898 181826 435454
rect 182382 434898 217826 435454
rect 218382 434898 253826 435454
rect 254382 434898 289826 435454
rect 290382 434898 325826 435454
rect 326382 434898 361826 435454
rect 362382 434898 397826 435454
rect 398382 434898 433826 435454
rect 434382 434898 469826 435454
rect 470382 434898 505826 435454
rect 506382 434898 541826 435454
rect 542382 434898 577826 435454
rect 578382 434898 585342 435454
rect 585898 434898 592650 435454
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 424938 -8694 425494
rect -8138 424938 27866 425494
rect 28422 424938 63866 425494
rect 64422 424938 99866 425494
rect 100422 424938 135866 425494
rect 136422 424938 171866 425494
rect 172422 424938 207866 425494
rect 208422 424938 243866 425494
rect 244422 424938 279866 425494
rect 280422 424938 315866 425494
rect 316422 424938 351866 425494
rect 352422 424938 387866 425494
rect 388422 424938 423866 425494
rect 424422 424938 459866 425494
rect 460422 424938 495866 425494
rect 496422 424938 531866 425494
rect 532422 424938 567866 425494
rect 568422 424938 592062 425494
rect 592618 424938 592650 425494
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421218 -7734 421774
rect -7178 421218 24146 421774
rect 24702 421218 60146 421774
rect 60702 421218 96146 421774
rect 96702 421218 132146 421774
rect 132702 421218 168146 421774
rect 168702 421218 204146 421774
rect 204702 421218 240146 421774
rect 240702 421218 276146 421774
rect 276702 421218 312146 421774
rect 312702 421218 348146 421774
rect 348702 421218 384146 421774
rect 384702 421218 420146 421774
rect 420702 421218 456146 421774
rect 456702 421218 492146 421774
rect 492702 421218 528146 421774
rect 528702 421218 564146 421774
rect 564702 421218 591102 421774
rect 591658 421218 592650 421774
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417498 -6774 418054
rect -6218 417498 20426 418054
rect 20982 417498 56426 418054
rect 56982 417498 92426 418054
rect 92982 417498 128426 418054
rect 128982 417498 164426 418054
rect 164982 417498 200426 418054
rect 200982 417498 236426 418054
rect 236982 417498 272426 418054
rect 272982 417498 308426 418054
rect 308982 417498 344426 418054
rect 344982 417498 380426 418054
rect 380982 417498 416426 418054
rect 416982 417498 452426 418054
rect 452982 417498 488426 418054
rect 488982 417498 524426 418054
rect 524982 417498 560426 418054
rect 560982 417498 590142 418054
rect 590698 417498 592650 418054
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 413778 -5814 414334
rect -5258 413778 16706 414334
rect 17262 413778 52706 414334
rect 53262 413778 88706 414334
rect 89262 413778 124706 414334
rect 125262 413778 160706 414334
rect 161262 413778 196706 414334
rect 197262 413778 232706 414334
rect 233262 413778 268706 414334
rect 269262 413778 304706 414334
rect 305262 413778 340706 414334
rect 341262 413778 376706 414334
rect 377262 413778 412706 414334
rect 413262 413778 448706 414334
rect 449262 413778 484706 414334
rect 485262 413778 520706 414334
rect 521262 413778 556706 414334
rect 557262 413778 589182 414334
rect 589738 413778 592650 414334
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410058 -4854 410614
rect -4298 410058 12986 410614
rect 13542 410058 48986 410614
rect 49542 410058 84986 410614
rect 85542 410058 120986 410614
rect 121542 410058 156986 410614
rect 157542 410058 192986 410614
rect 193542 410058 228986 410614
rect 229542 410058 264986 410614
rect 265542 410058 300986 410614
rect 301542 410058 336986 410614
rect 337542 410058 372986 410614
rect 373542 410058 408986 410614
rect 409542 410058 444986 410614
rect 445542 410058 480986 410614
rect 481542 410058 516986 410614
rect 517542 410058 552986 410614
rect 553542 410058 588222 410614
rect 588778 410058 592650 410614
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406338 -3894 406894
rect -3338 406338 9266 406894
rect 9822 406338 45266 406894
rect 45822 406338 81266 406894
rect 81822 406338 117266 406894
rect 117822 406338 153266 406894
rect 153822 406338 189266 406894
rect 189822 406338 225266 406894
rect 225822 406338 261266 406894
rect 261822 406338 297266 406894
rect 297822 406338 333266 406894
rect 333822 406338 369266 406894
rect 369822 406338 405266 406894
rect 405822 406338 441266 406894
rect 441822 406338 477266 406894
rect 477822 406338 513266 406894
rect 513822 406338 549266 406894
rect 549822 406338 587262 406894
rect 587818 406338 592650 406894
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402618 -2934 403174
rect -2378 402618 5546 403174
rect 6102 402618 41546 403174
rect 42102 402618 77546 403174
rect 78102 402618 113546 403174
rect 114102 402618 149546 403174
rect 150102 402618 185546 403174
rect 186102 402618 221546 403174
rect 222102 402618 257546 403174
rect 258102 402618 293546 403174
rect 294102 402618 329546 403174
rect 330102 402618 365546 403174
rect 366102 402618 401546 403174
rect 402102 402618 437546 403174
rect 438102 402618 473546 403174
rect 474102 402618 509546 403174
rect 510102 402618 545546 403174
rect 546102 402618 581546 403174
rect 582102 402618 586302 403174
rect 586858 402618 592650 403174
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 398898 -1974 399454
rect -1418 398898 1826 399454
rect 2382 398898 37826 399454
rect 38382 398898 73826 399454
rect 74382 398898 109826 399454
rect 110382 398898 145826 399454
rect 146382 398898 181826 399454
rect 182382 398898 217826 399454
rect 218382 398898 253826 399454
rect 254382 398898 289826 399454
rect 290382 398898 325826 399454
rect 326382 398898 361826 399454
rect 362382 398898 397826 399454
rect 398382 398898 433826 399454
rect 434382 398898 469826 399454
rect 470382 398898 505826 399454
rect 506382 398898 541826 399454
rect 542382 398898 577826 399454
rect 578382 398898 585342 399454
rect 585898 398898 592650 399454
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 388938 -8694 389494
rect -8138 388938 27866 389494
rect 28422 388938 63866 389494
rect 64422 388938 99866 389494
rect 100422 388938 135866 389494
rect 136422 388938 171866 389494
rect 172422 388938 207866 389494
rect 208422 388938 243866 389494
rect 244422 388938 279866 389494
rect 280422 388938 315866 389494
rect 316422 388938 351866 389494
rect 352422 388938 387866 389494
rect 388422 388938 423866 389494
rect 424422 388938 459866 389494
rect 460422 388938 495866 389494
rect 496422 388938 531866 389494
rect 532422 388938 567866 389494
rect 568422 388938 592062 389494
rect 592618 388938 592650 389494
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385218 -7734 385774
rect -7178 385218 24146 385774
rect 24702 385218 60146 385774
rect 60702 385218 96146 385774
rect 96702 385218 132146 385774
rect 132702 385218 168146 385774
rect 168702 385218 204146 385774
rect 204702 385218 240146 385774
rect 240702 385218 276146 385774
rect 276702 385218 312146 385774
rect 312702 385218 348146 385774
rect 348702 385218 384146 385774
rect 384702 385218 420146 385774
rect 420702 385218 456146 385774
rect 456702 385218 492146 385774
rect 492702 385218 528146 385774
rect 528702 385218 564146 385774
rect 564702 385218 591102 385774
rect 591658 385218 592650 385774
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381498 -6774 382054
rect -6218 381498 20426 382054
rect 20982 381498 56426 382054
rect 56982 381498 92426 382054
rect 92982 381498 128426 382054
rect 128982 381498 164426 382054
rect 164982 381498 200426 382054
rect 200982 381498 236426 382054
rect 236982 381498 272426 382054
rect 272982 381498 308426 382054
rect 308982 381498 344426 382054
rect 344982 381498 380426 382054
rect 380982 381498 416426 382054
rect 416982 381498 452426 382054
rect 452982 381498 488426 382054
rect 488982 381498 524426 382054
rect 524982 381498 560426 382054
rect 560982 381498 590142 382054
rect 590698 381498 592650 382054
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 377778 -5814 378334
rect -5258 377778 16706 378334
rect 17262 377778 52706 378334
rect 53262 377778 88706 378334
rect 89262 377778 124706 378334
rect 125262 377778 160706 378334
rect 161262 377778 196706 378334
rect 197262 377778 232706 378334
rect 233262 377778 268706 378334
rect 269262 377778 304706 378334
rect 305262 377778 340706 378334
rect 341262 377778 376706 378334
rect 377262 377778 412706 378334
rect 413262 377778 448706 378334
rect 449262 377778 484706 378334
rect 485262 377778 520706 378334
rect 521262 377778 556706 378334
rect 557262 377778 589182 378334
rect 589738 377778 592650 378334
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374058 -4854 374614
rect -4298 374058 12986 374614
rect 13542 374058 48986 374614
rect 49542 374058 84986 374614
rect 85542 374058 120986 374614
rect 121542 374058 156986 374614
rect 157542 374058 192986 374614
rect 193542 374058 228986 374614
rect 229542 374058 264986 374614
rect 265542 374058 300986 374614
rect 301542 374058 336986 374614
rect 337542 374058 372986 374614
rect 373542 374058 408986 374614
rect 409542 374058 444986 374614
rect 445542 374058 480986 374614
rect 481542 374058 516986 374614
rect 517542 374058 552986 374614
rect 553542 374058 588222 374614
rect 588778 374058 592650 374614
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370338 -3894 370894
rect -3338 370338 9266 370894
rect 9822 370338 45266 370894
rect 45822 370338 81266 370894
rect 81822 370338 117266 370894
rect 117822 370338 153266 370894
rect 153822 370338 189266 370894
rect 189822 370338 225266 370894
rect 225822 370338 261266 370894
rect 261822 370338 297266 370894
rect 297822 370338 333266 370894
rect 333822 370338 369266 370894
rect 369822 370338 405266 370894
rect 405822 370338 441266 370894
rect 441822 370338 477266 370894
rect 477822 370338 513266 370894
rect 513822 370338 549266 370894
rect 549822 370338 587262 370894
rect 587818 370338 592650 370894
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366618 -2934 367174
rect -2378 366618 5546 367174
rect 6102 366618 41546 367174
rect 42102 366618 77546 367174
rect 78102 366618 113546 367174
rect 114102 366618 149546 367174
rect 150102 366618 185546 367174
rect 186102 366618 221546 367174
rect 222102 366618 257546 367174
rect 258102 366618 293546 367174
rect 294102 366618 329546 367174
rect 330102 366618 365546 367174
rect 366102 366618 401546 367174
rect 402102 366618 437546 367174
rect 438102 366618 473546 367174
rect 474102 366618 509546 367174
rect 510102 366618 545546 367174
rect 546102 366618 581546 367174
rect 582102 366618 586302 367174
rect 586858 366618 592650 367174
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 362898 -1974 363454
rect -1418 362898 1826 363454
rect 2382 362898 37826 363454
rect 38382 362898 73826 363454
rect 74382 362898 109826 363454
rect 110382 362898 145826 363454
rect 146382 362898 181826 363454
rect 182382 362898 217826 363454
rect 218382 362898 253826 363454
rect 254382 362898 289826 363454
rect 290382 362898 325826 363454
rect 326382 362898 361826 363454
rect 362382 362898 397826 363454
rect 398382 362898 433826 363454
rect 434382 362898 469826 363454
rect 470382 362898 505826 363454
rect 506382 362898 541826 363454
rect 542382 362898 577826 363454
rect 578382 362898 585342 363454
rect 585898 362898 592650 363454
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 352938 -8694 353494
rect -8138 352938 27866 353494
rect 28422 352938 63866 353494
rect 64422 352938 99866 353494
rect 100422 352938 135866 353494
rect 136422 352938 171866 353494
rect 172422 352938 207866 353494
rect 208422 352938 243866 353494
rect 244422 352938 279866 353494
rect 280422 352938 315866 353494
rect 316422 352938 351866 353494
rect 352422 352938 387866 353494
rect 388422 352938 423866 353494
rect 424422 352938 459866 353494
rect 460422 352938 495866 353494
rect 496422 352938 531866 353494
rect 532422 352938 567866 353494
rect 568422 352938 592062 353494
rect 592618 352938 592650 353494
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349218 -7734 349774
rect -7178 349218 24146 349774
rect 24702 349218 60146 349774
rect 60702 349218 96146 349774
rect 96702 349218 132146 349774
rect 132702 349218 168146 349774
rect 168702 349218 204146 349774
rect 204702 349218 240146 349774
rect 240702 349218 276146 349774
rect 276702 349218 312146 349774
rect 312702 349218 348146 349774
rect 348702 349218 420146 349774
rect 420702 349218 456146 349774
rect 456702 349218 528146 349774
rect 528702 349218 564146 349774
rect 564702 349218 591102 349774
rect 591658 349218 592650 349774
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345498 -6774 346054
rect -6218 345498 20426 346054
rect 20982 345498 56426 346054
rect 56982 345498 128426 346054
rect 128982 345498 164426 346054
rect 164982 345498 236426 346054
rect 236982 345498 272426 346054
rect 272982 345498 344426 346054
rect 344982 345498 380426 346054
rect 380982 345498 416426 346054
rect 416982 345498 452426 346054
rect 452982 345498 488426 346054
rect 488982 345498 524426 346054
rect 524982 345498 560426 346054
rect 560982 345498 590142 346054
rect 590698 345498 592650 346054
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 341778 -5814 342334
rect -5258 341778 16706 342334
rect 17262 341778 52706 342334
rect 53262 341778 88706 342334
rect 89262 341778 124706 342334
rect 125262 341778 160706 342334
rect 161262 341778 196706 342334
rect 197262 341778 232706 342334
rect 233262 341778 268706 342334
rect 269262 341778 304706 342334
rect 305262 341778 340706 342334
rect 341262 341778 376706 342334
rect 377262 341778 412706 342334
rect 413262 341778 448706 342334
rect 449262 341778 484706 342334
rect 485262 341778 520706 342334
rect 521262 341778 556706 342334
rect 557262 341778 589182 342334
rect 589738 341778 592650 342334
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338058 -4854 338614
rect -4298 338058 12986 338614
rect 13542 338058 48986 338614
rect 49542 338058 84986 338614
rect 85542 338058 120986 338614
rect 121542 338058 156986 338614
rect 157542 338058 192986 338614
rect 193542 338058 228986 338614
rect 229542 338058 264986 338614
rect 265542 338058 300986 338614
rect 301542 338058 336986 338614
rect 337542 338058 372986 338614
rect 373542 338058 408986 338614
rect 409542 338058 444986 338614
rect 445542 338058 480986 338614
rect 481542 338058 516986 338614
rect 517542 338058 552986 338614
rect 553542 338058 588222 338614
rect 588778 338058 592650 338614
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334338 -3894 334894
rect -3338 334338 9266 334894
rect 9822 334338 45266 334894
rect 45822 334338 81266 334894
rect 81822 334338 117266 334894
rect 117822 334338 153266 334894
rect 153822 334338 189266 334894
rect 189822 334338 225266 334894
rect 225822 334338 297266 334894
rect 297822 334338 333266 334894
rect 333822 334338 405266 334894
rect 405822 334338 441266 334894
rect 441822 334338 513266 334894
rect 513822 334338 549266 334894
rect 549822 334338 587262 334894
rect 587818 334338 592650 334894
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330618 -2934 331174
rect -2378 330618 5546 331174
rect 6102 330938 31610 331174
rect 31846 330938 41546 331174
rect 6102 330854 41546 330938
rect 6102 330618 31610 330854
rect 31846 330618 41546 330854
rect 42102 330938 62330 331174
rect 62566 330938 93050 331174
rect 93286 330938 113546 331174
rect 42102 330854 113546 330938
rect 42102 330618 62330 330854
rect 62566 330618 93050 330854
rect 93286 330618 113546 330854
rect 114102 330938 123770 331174
rect 124006 330938 149546 331174
rect 114102 330854 149546 330938
rect 114102 330618 123770 330854
rect 124006 330618 149546 330854
rect 150102 330938 154490 331174
rect 154726 330938 185210 331174
rect 185446 330938 215930 331174
rect 216166 330938 221546 331174
rect 150102 330854 221546 330938
rect 150102 330618 154490 330854
rect 154726 330618 185210 330854
rect 185446 330618 215930 330854
rect 216166 330618 221546 330854
rect 222102 330938 246650 331174
rect 246886 330938 257546 331174
rect 222102 330854 257546 330938
rect 222102 330618 246650 330854
rect 246886 330618 257546 330854
rect 258102 330938 277370 331174
rect 277606 330938 293546 331174
rect 258102 330854 293546 330938
rect 258102 330618 277370 330854
rect 277606 330618 293546 330854
rect 294102 330938 308090 331174
rect 308326 330938 329546 331174
rect 294102 330854 329546 330938
rect 294102 330618 308090 330854
rect 308326 330618 329546 330854
rect 330102 330938 338810 331174
rect 339046 330938 365546 331174
rect 330102 330854 365546 330938
rect 330102 330618 338810 330854
rect 339046 330618 365546 330854
rect 366102 330938 369530 331174
rect 369766 330938 400250 331174
rect 400486 330938 401546 331174
rect 366102 330854 401546 330938
rect 366102 330618 369530 330854
rect 369766 330618 400250 330854
rect 400486 330618 401546 330854
rect 402102 330938 430970 331174
rect 431206 330938 437546 331174
rect 402102 330854 437546 330938
rect 402102 330618 430970 330854
rect 431206 330618 437546 330854
rect 438102 330938 461690 331174
rect 461926 330938 473546 331174
rect 438102 330854 473546 330938
rect 438102 330618 461690 330854
rect 461926 330618 473546 330854
rect 474102 330938 492410 331174
rect 492646 330938 509546 331174
rect 474102 330854 509546 330938
rect 474102 330618 492410 330854
rect 492646 330618 509546 330854
rect 510102 330938 523130 331174
rect 523366 330938 545546 331174
rect 510102 330854 545546 330938
rect 510102 330618 523130 330854
rect 523366 330618 545546 330854
rect 546102 330938 553850 331174
rect 554086 330938 581546 331174
rect 546102 330854 581546 330938
rect 546102 330618 553850 330854
rect 554086 330618 581546 330854
rect 582102 330618 586302 331174
rect 586858 330618 592650 331174
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 326898 -1974 327454
rect -1418 326898 1826 327454
rect 2382 327218 16250 327454
rect 16486 327218 37826 327454
rect 2382 327134 37826 327218
rect 2382 326898 16250 327134
rect 16486 326898 37826 327134
rect 38382 327218 46970 327454
rect 47206 327218 73826 327454
rect 38382 327134 73826 327218
rect 38382 326898 46970 327134
rect 47206 326898 73826 327134
rect 74382 327218 77690 327454
rect 77926 327218 108410 327454
rect 108646 327218 109826 327454
rect 74382 327134 109826 327218
rect 74382 326898 77690 327134
rect 77926 326898 108410 327134
rect 108646 326898 109826 327134
rect 110382 327218 139130 327454
rect 139366 327218 145826 327454
rect 110382 327134 145826 327218
rect 110382 326898 139130 327134
rect 139366 326898 145826 327134
rect 146382 327218 169850 327454
rect 170086 327218 181826 327454
rect 146382 327134 181826 327218
rect 146382 326898 169850 327134
rect 170086 326898 181826 327134
rect 182382 327218 200570 327454
rect 200806 327218 217826 327454
rect 182382 327134 217826 327218
rect 182382 326898 200570 327134
rect 200806 326898 217826 327134
rect 218382 327218 231290 327454
rect 231526 327218 253826 327454
rect 218382 327134 253826 327218
rect 218382 326898 231290 327134
rect 231526 326898 253826 327134
rect 254382 327218 262010 327454
rect 262246 327218 289826 327454
rect 254382 327134 289826 327218
rect 254382 326898 262010 327134
rect 262246 326898 289826 327134
rect 290382 327218 292730 327454
rect 292966 327218 323450 327454
rect 323686 327218 325826 327454
rect 290382 327134 325826 327218
rect 290382 326898 292730 327134
rect 292966 326898 323450 327134
rect 323686 326898 325826 327134
rect 326382 327218 354170 327454
rect 354406 327218 361826 327454
rect 326382 327134 361826 327218
rect 326382 326898 354170 327134
rect 354406 326898 361826 327134
rect 362382 327218 384890 327454
rect 385126 327218 397826 327454
rect 362382 327134 397826 327218
rect 362382 326898 384890 327134
rect 385126 326898 397826 327134
rect 398382 327218 415610 327454
rect 415846 327218 433826 327454
rect 398382 327134 433826 327218
rect 398382 326898 415610 327134
rect 415846 326898 433826 327134
rect 434382 327218 446330 327454
rect 446566 327218 469826 327454
rect 434382 327134 469826 327218
rect 434382 326898 446330 327134
rect 446566 326898 469826 327134
rect 470382 327218 477050 327454
rect 477286 327218 505826 327454
rect 470382 327134 505826 327218
rect 470382 326898 477050 327134
rect 477286 326898 505826 327134
rect 506382 327218 507770 327454
rect 508006 327218 538490 327454
rect 538726 327218 541826 327454
rect 506382 327134 541826 327218
rect 506382 326898 507770 327134
rect 508006 326898 538490 327134
rect 538726 326898 541826 327134
rect 542382 327218 569210 327454
rect 569446 327218 577826 327454
rect 542382 327134 577826 327218
rect 542382 326898 569210 327134
rect 569446 326898 577826 327134
rect 578382 326898 585342 327454
rect 585898 326898 592650 327454
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 316938 -8694 317494
rect -8138 316938 27866 317494
rect 28422 316938 63866 317494
rect 64422 316938 99866 317494
rect 100422 316938 135866 317494
rect 136422 316938 171866 317494
rect 172422 316938 207866 317494
rect 208422 316938 243866 317494
rect 244422 316938 279866 317494
rect 280422 316938 315866 317494
rect 316422 316938 351866 317494
rect 352422 316938 387866 317494
rect 388422 316938 423866 317494
rect 424422 316938 459866 317494
rect 460422 316938 495866 317494
rect 496422 316938 531866 317494
rect 532422 316938 567866 317494
rect 568422 316938 592062 317494
rect 592618 316938 592650 317494
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313218 -7734 313774
rect -7178 313218 24146 313774
rect 24702 313218 60146 313774
rect 60702 313218 96146 313774
rect 96702 313218 132146 313774
rect 132702 313218 168146 313774
rect 168702 313218 204146 313774
rect 204702 313218 240146 313774
rect 240702 313218 276146 313774
rect 276702 313218 312146 313774
rect 312702 313218 348146 313774
rect 348702 313218 420146 313774
rect 420702 313218 456146 313774
rect 456702 313218 528146 313774
rect 528702 313218 564146 313774
rect 564702 313218 591102 313774
rect 591658 313218 592650 313774
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309498 -6774 310054
rect -6218 309498 20426 310054
rect 20982 309498 56426 310054
rect 56982 309498 128426 310054
rect 128982 309498 164426 310054
rect 164982 309498 236426 310054
rect 236982 309498 272426 310054
rect 272982 309498 344426 310054
rect 344982 309498 380426 310054
rect 380982 309498 416426 310054
rect 416982 309498 452426 310054
rect 452982 309498 488426 310054
rect 488982 309498 524426 310054
rect 524982 309498 560426 310054
rect 560982 309498 590142 310054
rect 590698 309498 592650 310054
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 305778 -5814 306334
rect -5258 305778 16706 306334
rect 17262 305778 52706 306334
rect 53262 305778 88706 306334
rect 89262 305778 124706 306334
rect 125262 305778 160706 306334
rect 161262 305778 196706 306334
rect 197262 305778 232706 306334
rect 233262 305778 268706 306334
rect 269262 305778 304706 306334
rect 305262 305778 340706 306334
rect 341262 305778 376706 306334
rect 377262 305778 412706 306334
rect 413262 305778 448706 306334
rect 449262 305778 484706 306334
rect 485262 305778 520706 306334
rect 521262 305778 556706 306334
rect 557262 305778 589182 306334
rect 589738 305778 592650 306334
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302058 -4854 302614
rect -4298 302058 12986 302614
rect 13542 302058 48986 302614
rect 49542 302058 84986 302614
rect 85542 302058 120986 302614
rect 121542 302058 156986 302614
rect 157542 302058 192986 302614
rect 193542 302058 228986 302614
rect 229542 302058 264986 302614
rect 265542 302058 300986 302614
rect 301542 302058 336986 302614
rect 337542 302058 372986 302614
rect 373542 302058 408986 302614
rect 409542 302058 444986 302614
rect 445542 302058 480986 302614
rect 481542 302058 516986 302614
rect 517542 302058 552986 302614
rect 553542 302058 588222 302614
rect 588778 302058 592650 302614
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298338 -3894 298894
rect -3338 298338 9266 298894
rect 9822 298338 45266 298894
rect 45822 298338 81266 298894
rect 81822 298338 117266 298894
rect 117822 298338 153266 298894
rect 153822 298338 189266 298894
rect 189822 298338 225266 298894
rect 225822 298338 297266 298894
rect 297822 298338 333266 298894
rect 333822 298338 405266 298894
rect 405822 298338 441266 298894
rect 441822 298338 513266 298894
rect 513822 298338 549266 298894
rect 549822 298338 587262 298894
rect 587818 298338 592650 298894
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294618 -2934 295174
rect -2378 294618 5546 295174
rect 6102 294938 31610 295174
rect 31846 294938 41546 295174
rect 6102 294854 41546 294938
rect 6102 294618 31610 294854
rect 31846 294618 41546 294854
rect 42102 294938 62330 295174
rect 62566 294938 93050 295174
rect 93286 294938 113546 295174
rect 42102 294854 113546 294938
rect 42102 294618 62330 294854
rect 62566 294618 93050 294854
rect 93286 294618 113546 294854
rect 114102 294938 123770 295174
rect 124006 294938 149546 295174
rect 114102 294854 149546 294938
rect 114102 294618 123770 294854
rect 124006 294618 149546 294854
rect 150102 294938 154490 295174
rect 154726 294938 185210 295174
rect 185446 294938 215930 295174
rect 216166 294938 221546 295174
rect 150102 294854 221546 294938
rect 150102 294618 154490 294854
rect 154726 294618 185210 294854
rect 185446 294618 215930 294854
rect 216166 294618 221546 294854
rect 222102 294938 246650 295174
rect 246886 294938 257546 295174
rect 222102 294854 257546 294938
rect 222102 294618 246650 294854
rect 246886 294618 257546 294854
rect 258102 294938 277370 295174
rect 277606 294938 293546 295174
rect 258102 294854 293546 294938
rect 258102 294618 277370 294854
rect 277606 294618 293546 294854
rect 294102 294938 308090 295174
rect 308326 294938 329546 295174
rect 294102 294854 329546 294938
rect 294102 294618 308090 294854
rect 308326 294618 329546 294854
rect 330102 294938 338810 295174
rect 339046 294938 365546 295174
rect 330102 294854 365546 294938
rect 330102 294618 338810 294854
rect 339046 294618 365546 294854
rect 366102 294938 369530 295174
rect 369766 294938 400250 295174
rect 400486 294938 401546 295174
rect 366102 294854 401546 294938
rect 366102 294618 369530 294854
rect 369766 294618 400250 294854
rect 400486 294618 401546 294854
rect 402102 294938 430970 295174
rect 431206 294938 437546 295174
rect 402102 294854 437546 294938
rect 402102 294618 430970 294854
rect 431206 294618 437546 294854
rect 438102 294938 461690 295174
rect 461926 294938 473546 295174
rect 438102 294854 473546 294938
rect 438102 294618 461690 294854
rect 461926 294618 473546 294854
rect 474102 294938 492410 295174
rect 492646 294938 509546 295174
rect 474102 294854 509546 294938
rect 474102 294618 492410 294854
rect 492646 294618 509546 294854
rect 510102 294938 523130 295174
rect 523366 294938 545546 295174
rect 510102 294854 545546 294938
rect 510102 294618 523130 294854
rect 523366 294618 545546 294854
rect 546102 294938 553850 295174
rect 554086 294938 581546 295174
rect 546102 294854 581546 294938
rect 546102 294618 553850 294854
rect 554086 294618 581546 294854
rect 582102 294618 586302 295174
rect 586858 294618 592650 295174
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 290898 -1974 291454
rect -1418 290898 1826 291454
rect 2382 291218 16250 291454
rect 16486 291218 37826 291454
rect 2382 291134 37826 291218
rect 2382 290898 16250 291134
rect 16486 290898 37826 291134
rect 38382 291218 46970 291454
rect 47206 291218 73826 291454
rect 38382 291134 73826 291218
rect 38382 290898 46970 291134
rect 47206 290898 73826 291134
rect 74382 291218 77690 291454
rect 77926 291218 108410 291454
rect 108646 291218 109826 291454
rect 74382 291134 109826 291218
rect 74382 290898 77690 291134
rect 77926 290898 108410 291134
rect 108646 290898 109826 291134
rect 110382 291218 139130 291454
rect 139366 291218 145826 291454
rect 110382 291134 145826 291218
rect 110382 290898 139130 291134
rect 139366 290898 145826 291134
rect 146382 291218 169850 291454
rect 170086 291218 181826 291454
rect 146382 291134 181826 291218
rect 146382 290898 169850 291134
rect 170086 290898 181826 291134
rect 182382 291218 200570 291454
rect 200806 291218 217826 291454
rect 182382 291134 217826 291218
rect 182382 290898 200570 291134
rect 200806 290898 217826 291134
rect 218382 291218 231290 291454
rect 231526 291218 253826 291454
rect 218382 291134 253826 291218
rect 218382 290898 231290 291134
rect 231526 290898 253826 291134
rect 254382 291218 262010 291454
rect 262246 291218 289826 291454
rect 254382 291134 289826 291218
rect 254382 290898 262010 291134
rect 262246 290898 289826 291134
rect 290382 291218 292730 291454
rect 292966 291218 323450 291454
rect 323686 291218 325826 291454
rect 290382 291134 325826 291218
rect 290382 290898 292730 291134
rect 292966 290898 323450 291134
rect 323686 290898 325826 291134
rect 326382 291218 354170 291454
rect 354406 291218 361826 291454
rect 326382 291134 361826 291218
rect 326382 290898 354170 291134
rect 354406 290898 361826 291134
rect 362382 291218 384890 291454
rect 385126 291218 397826 291454
rect 362382 291134 397826 291218
rect 362382 290898 384890 291134
rect 385126 290898 397826 291134
rect 398382 291218 415610 291454
rect 415846 291218 433826 291454
rect 398382 291134 433826 291218
rect 398382 290898 415610 291134
rect 415846 290898 433826 291134
rect 434382 291218 446330 291454
rect 446566 291218 469826 291454
rect 434382 291134 469826 291218
rect 434382 290898 446330 291134
rect 446566 290898 469826 291134
rect 470382 291218 477050 291454
rect 477286 291218 505826 291454
rect 470382 291134 505826 291218
rect 470382 290898 477050 291134
rect 477286 290898 505826 291134
rect 506382 291218 507770 291454
rect 508006 291218 538490 291454
rect 538726 291218 541826 291454
rect 506382 291134 541826 291218
rect 506382 290898 507770 291134
rect 508006 290898 538490 291134
rect 538726 290898 541826 291134
rect 542382 291218 569210 291454
rect 569446 291218 577826 291454
rect 542382 291134 577826 291218
rect 542382 290898 569210 291134
rect 569446 290898 577826 291134
rect 578382 290898 585342 291454
rect 585898 290898 592650 291454
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 280938 -8694 281494
rect -8138 280938 27866 281494
rect 28422 280938 63866 281494
rect 64422 280938 99866 281494
rect 100422 280938 135866 281494
rect 136422 280938 171866 281494
rect 172422 280938 207866 281494
rect 208422 280938 243866 281494
rect 244422 280938 279866 281494
rect 280422 280938 315866 281494
rect 316422 280938 351866 281494
rect 352422 280938 387866 281494
rect 388422 280938 423866 281494
rect 424422 280938 459866 281494
rect 460422 280938 495866 281494
rect 496422 280938 531866 281494
rect 532422 280938 567866 281494
rect 568422 280938 592062 281494
rect 592618 280938 592650 281494
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277218 -7734 277774
rect -7178 277218 24146 277774
rect 24702 277218 60146 277774
rect 60702 277218 96146 277774
rect 96702 277218 132146 277774
rect 132702 277218 168146 277774
rect 168702 277218 204146 277774
rect 204702 277218 240146 277774
rect 240702 277218 276146 277774
rect 276702 277218 312146 277774
rect 312702 277218 348146 277774
rect 348702 277218 420146 277774
rect 420702 277218 456146 277774
rect 456702 277218 528146 277774
rect 528702 277218 564146 277774
rect 564702 277218 591102 277774
rect 591658 277218 592650 277774
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273498 -6774 274054
rect -6218 273498 20426 274054
rect 20982 273498 56426 274054
rect 56982 273498 128426 274054
rect 128982 273498 164426 274054
rect 164982 273498 236426 274054
rect 236982 273498 272426 274054
rect 272982 273498 344426 274054
rect 344982 273498 380426 274054
rect 380982 273498 416426 274054
rect 416982 273498 452426 274054
rect 452982 273498 488426 274054
rect 488982 273498 524426 274054
rect 524982 273498 560426 274054
rect 560982 273498 590142 274054
rect 590698 273498 592650 274054
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 269778 -5814 270334
rect -5258 269778 16706 270334
rect 17262 269778 52706 270334
rect 53262 269778 88706 270334
rect 89262 269778 124706 270334
rect 125262 269778 160706 270334
rect 161262 269778 196706 270334
rect 197262 269778 232706 270334
rect 233262 269778 268706 270334
rect 269262 269778 304706 270334
rect 305262 269778 340706 270334
rect 341262 269778 376706 270334
rect 377262 269778 412706 270334
rect 413262 269778 448706 270334
rect 449262 269778 484706 270334
rect 485262 269778 520706 270334
rect 521262 269778 556706 270334
rect 557262 269778 589182 270334
rect 589738 269778 592650 270334
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266058 -4854 266614
rect -4298 266058 12986 266614
rect 13542 266058 48986 266614
rect 49542 266058 84986 266614
rect 85542 266058 120986 266614
rect 121542 266058 156986 266614
rect 157542 266058 192986 266614
rect 193542 266058 228986 266614
rect 229542 266058 264986 266614
rect 265542 266058 300986 266614
rect 301542 266058 336986 266614
rect 337542 266058 372986 266614
rect 373542 266058 408986 266614
rect 409542 266058 444986 266614
rect 445542 266058 480986 266614
rect 481542 266058 516986 266614
rect 517542 266058 552986 266614
rect 553542 266058 588222 266614
rect 588778 266058 592650 266614
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262338 -3894 262894
rect -3338 262338 9266 262894
rect 9822 262338 45266 262894
rect 45822 262338 81266 262894
rect 81822 262338 117266 262894
rect 117822 262338 153266 262894
rect 153822 262338 189266 262894
rect 189822 262338 225266 262894
rect 225822 262338 297266 262894
rect 297822 262338 333266 262894
rect 333822 262338 405266 262894
rect 405822 262338 441266 262894
rect 441822 262338 513266 262894
rect 513822 262338 549266 262894
rect 549822 262338 587262 262894
rect 587818 262338 592650 262894
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258618 -2934 259174
rect -2378 258618 5546 259174
rect 6102 258938 31610 259174
rect 31846 258938 41546 259174
rect 6102 258854 41546 258938
rect 6102 258618 31610 258854
rect 31846 258618 41546 258854
rect 42102 258938 62330 259174
rect 62566 258938 93050 259174
rect 93286 258938 113546 259174
rect 42102 258854 113546 258938
rect 42102 258618 62330 258854
rect 62566 258618 93050 258854
rect 93286 258618 113546 258854
rect 114102 258938 123770 259174
rect 124006 258938 149546 259174
rect 114102 258854 149546 258938
rect 114102 258618 123770 258854
rect 124006 258618 149546 258854
rect 150102 258938 154490 259174
rect 154726 258938 185210 259174
rect 185446 258938 215930 259174
rect 216166 258938 221546 259174
rect 150102 258854 221546 258938
rect 150102 258618 154490 258854
rect 154726 258618 185210 258854
rect 185446 258618 215930 258854
rect 216166 258618 221546 258854
rect 222102 258938 246650 259174
rect 246886 258938 257546 259174
rect 222102 258854 257546 258938
rect 222102 258618 246650 258854
rect 246886 258618 257546 258854
rect 258102 258938 277370 259174
rect 277606 258938 293546 259174
rect 258102 258854 293546 258938
rect 258102 258618 277370 258854
rect 277606 258618 293546 258854
rect 294102 258938 308090 259174
rect 308326 258938 329546 259174
rect 294102 258854 329546 258938
rect 294102 258618 308090 258854
rect 308326 258618 329546 258854
rect 330102 258938 338810 259174
rect 339046 258938 365546 259174
rect 330102 258854 365546 258938
rect 330102 258618 338810 258854
rect 339046 258618 365546 258854
rect 366102 258938 369530 259174
rect 369766 258938 400250 259174
rect 400486 258938 401546 259174
rect 366102 258854 401546 258938
rect 366102 258618 369530 258854
rect 369766 258618 400250 258854
rect 400486 258618 401546 258854
rect 402102 258938 430970 259174
rect 431206 258938 437546 259174
rect 402102 258854 437546 258938
rect 402102 258618 430970 258854
rect 431206 258618 437546 258854
rect 438102 258938 461690 259174
rect 461926 258938 473546 259174
rect 438102 258854 473546 258938
rect 438102 258618 461690 258854
rect 461926 258618 473546 258854
rect 474102 258938 492410 259174
rect 492646 258938 509546 259174
rect 474102 258854 509546 258938
rect 474102 258618 492410 258854
rect 492646 258618 509546 258854
rect 510102 258938 523130 259174
rect 523366 258938 545546 259174
rect 510102 258854 545546 258938
rect 510102 258618 523130 258854
rect 523366 258618 545546 258854
rect 546102 258938 553850 259174
rect 554086 258938 581546 259174
rect 546102 258854 581546 258938
rect 546102 258618 553850 258854
rect 554086 258618 581546 258854
rect 582102 258618 586302 259174
rect 586858 258618 592650 259174
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 254898 -1974 255454
rect -1418 254898 1826 255454
rect 2382 255218 16250 255454
rect 16486 255218 37826 255454
rect 2382 255134 37826 255218
rect 2382 254898 16250 255134
rect 16486 254898 37826 255134
rect 38382 255218 46970 255454
rect 47206 255218 73826 255454
rect 38382 255134 73826 255218
rect 38382 254898 46970 255134
rect 47206 254898 73826 255134
rect 74382 255218 77690 255454
rect 77926 255218 108410 255454
rect 108646 255218 109826 255454
rect 74382 255134 109826 255218
rect 74382 254898 77690 255134
rect 77926 254898 108410 255134
rect 108646 254898 109826 255134
rect 110382 255218 139130 255454
rect 139366 255218 145826 255454
rect 110382 255134 145826 255218
rect 110382 254898 139130 255134
rect 139366 254898 145826 255134
rect 146382 255218 169850 255454
rect 170086 255218 181826 255454
rect 146382 255134 181826 255218
rect 146382 254898 169850 255134
rect 170086 254898 181826 255134
rect 182382 255218 200570 255454
rect 200806 255218 217826 255454
rect 182382 255134 217826 255218
rect 182382 254898 200570 255134
rect 200806 254898 217826 255134
rect 218382 255218 231290 255454
rect 231526 255218 253826 255454
rect 218382 255134 253826 255218
rect 218382 254898 231290 255134
rect 231526 254898 253826 255134
rect 254382 255218 262010 255454
rect 262246 255218 289826 255454
rect 254382 255134 289826 255218
rect 254382 254898 262010 255134
rect 262246 254898 289826 255134
rect 290382 255218 292730 255454
rect 292966 255218 323450 255454
rect 323686 255218 325826 255454
rect 290382 255134 325826 255218
rect 290382 254898 292730 255134
rect 292966 254898 323450 255134
rect 323686 254898 325826 255134
rect 326382 255218 354170 255454
rect 354406 255218 361826 255454
rect 326382 255134 361826 255218
rect 326382 254898 354170 255134
rect 354406 254898 361826 255134
rect 362382 255218 384890 255454
rect 385126 255218 397826 255454
rect 362382 255134 397826 255218
rect 362382 254898 384890 255134
rect 385126 254898 397826 255134
rect 398382 255218 415610 255454
rect 415846 255218 433826 255454
rect 398382 255134 433826 255218
rect 398382 254898 415610 255134
rect 415846 254898 433826 255134
rect 434382 255218 446330 255454
rect 446566 255218 469826 255454
rect 434382 255134 469826 255218
rect 434382 254898 446330 255134
rect 446566 254898 469826 255134
rect 470382 255218 477050 255454
rect 477286 255218 505826 255454
rect 470382 255134 505826 255218
rect 470382 254898 477050 255134
rect 477286 254898 505826 255134
rect 506382 255218 507770 255454
rect 508006 255218 538490 255454
rect 538726 255218 541826 255454
rect 506382 255134 541826 255218
rect 506382 254898 507770 255134
rect 508006 254898 538490 255134
rect 538726 254898 541826 255134
rect 542382 255218 569210 255454
rect 569446 255218 577826 255454
rect 542382 255134 577826 255218
rect 542382 254898 569210 255134
rect 569446 254898 577826 255134
rect 578382 254898 585342 255454
rect 585898 254898 592650 255454
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 244938 -8694 245494
rect -8138 244938 27866 245494
rect 28422 244938 63866 245494
rect 64422 244938 99866 245494
rect 100422 244938 135866 245494
rect 136422 244938 171866 245494
rect 172422 244938 207866 245494
rect 208422 244938 243866 245494
rect 244422 244938 279866 245494
rect 280422 244938 315866 245494
rect 316422 244938 351866 245494
rect 352422 244938 387866 245494
rect 388422 244938 423866 245494
rect 424422 244938 459866 245494
rect 460422 244938 495866 245494
rect 496422 244938 531866 245494
rect 532422 244938 567866 245494
rect 568422 244938 592062 245494
rect 592618 244938 592650 245494
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241218 -7734 241774
rect -7178 241218 24146 241774
rect 24702 241218 60146 241774
rect 60702 241218 96146 241774
rect 96702 241218 132146 241774
rect 132702 241218 168146 241774
rect 168702 241218 204146 241774
rect 204702 241218 240146 241774
rect 240702 241218 276146 241774
rect 276702 241218 312146 241774
rect 312702 241218 348146 241774
rect 348702 241218 420146 241774
rect 420702 241218 456146 241774
rect 456702 241218 528146 241774
rect 528702 241218 564146 241774
rect 564702 241218 591102 241774
rect 591658 241218 592650 241774
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237498 -6774 238054
rect -6218 237498 20426 238054
rect 20982 237498 56426 238054
rect 56982 237498 128426 238054
rect 128982 237498 164426 238054
rect 164982 237498 236426 238054
rect 236982 237498 272426 238054
rect 272982 237498 344426 238054
rect 344982 237498 380426 238054
rect 380982 237498 416426 238054
rect 416982 237498 452426 238054
rect 452982 237498 488426 238054
rect 488982 237498 524426 238054
rect 524982 237498 560426 238054
rect 560982 237498 590142 238054
rect 590698 237498 592650 238054
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 233778 -5814 234334
rect -5258 233778 16706 234334
rect 17262 233778 52706 234334
rect 53262 233778 88706 234334
rect 89262 233778 124706 234334
rect 125262 233778 160706 234334
rect 161262 233778 196706 234334
rect 197262 233778 232706 234334
rect 233262 233778 268706 234334
rect 269262 233778 304706 234334
rect 305262 233778 340706 234334
rect 341262 233778 376706 234334
rect 377262 233778 412706 234334
rect 413262 233778 448706 234334
rect 449262 233778 484706 234334
rect 485262 233778 520706 234334
rect 521262 233778 556706 234334
rect 557262 233778 589182 234334
rect 589738 233778 592650 234334
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230058 -4854 230614
rect -4298 230058 12986 230614
rect 13542 230058 48986 230614
rect 49542 230058 84986 230614
rect 85542 230058 120986 230614
rect 121542 230058 156986 230614
rect 157542 230058 192986 230614
rect 193542 230058 228986 230614
rect 229542 230058 264986 230614
rect 265542 230058 300986 230614
rect 301542 230058 336986 230614
rect 337542 230058 372986 230614
rect 373542 230058 408986 230614
rect 409542 230058 444986 230614
rect 445542 230058 480986 230614
rect 481542 230058 516986 230614
rect 517542 230058 552986 230614
rect 553542 230058 588222 230614
rect 588778 230058 592650 230614
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226338 -3894 226894
rect -3338 226338 9266 226894
rect 9822 226338 45266 226894
rect 45822 226338 81266 226894
rect 81822 226338 117266 226894
rect 117822 226338 153266 226894
rect 153822 226338 189266 226894
rect 189822 226338 225266 226894
rect 225822 226338 297266 226894
rect 297822 226338 333266 226894
rect 333822 226338 405266 226894
rect 405822 226338 441266 226894
rect 441822 226338 513266 226894
rect 513822 226338 549266 226894
rect 549822 226338 587262 226894
rect 587818 226338 592650 226894
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222618 -2934 223174
rect -2378 222618 5546 223174
rect 6102 222938 31610 223174
rect 31846 222938 41546 223174
rect 6102 222854 41546 222938
rect 6102 222618 31610 222854
rect 31846 222618 41546 222854
rect 42102 222938 62330 223174
rect 62566 222938 93050 223174
rect 93286 222938 113546 223174
rect 42102 222854 113546 222938
rect 42102 222618 62330 222854
rect 62566 222618 93050 222854
rect 93286 222618 113546 222854
rect 114102 222938 123770 223174
rect 124006 222938 149546 223174
rect 114102 222854 149546 222938
rect 114102 222618 123770 222854
rect 124006 222618 149546 222854
rect 150102 222938 154490 223174
rect 154726 222938 185210 223174
rect 185446 222938 215930 223174
rect 216166 222938 221546 223174
rect 150102 222854 221546 222938
rect 150102 222618 154490 222854
rect 154726 222618 185210 222854
rect 185446 222618 215930 222854
rect 216166 222618 221546 222854
rect 222102 222938 246650 223174
rect 246886 222938 257546 223174
rect 222102 222854 257546 222938
rect 222102 222618 246650 222854
rect 246886 222618 257546 222854
rect 258102 222938 277370 223174
rect 277606 222938 293546 223174
rect 258102 222854 293546 222938
rect 258102 222618 277370 222854
rect 277606 222618 293546 222854
rect 294102 222938 308090 223174
rect 308326 222938 329546 223174
rect 294102 222854 329546 222938
rect 294102 222618 308090 222854
rect 308326 222618 329546 222854
rect 330102 222938 338810 223174
rect 339046 222938 365546 223174
rect 330102 222854 365546 222938
rect 330102 222618 338810 222854
rect 339046 222618 365546 222854
rect 366102 222938 369530 223174
rect 369766 222938 400250 223174
rect 400486 222938 401546 223174
rect 366102 222854 401546 222938
rect 366102 222618 369530 222854
rect 369766 222618 400250 222854
rect 400486 222618 401546 222854
rect 402102 222938 430970 223174
rect 431206 222938 437546 223174
rect 402102 222854 437546 222938
rect 402102 222618 430970 222854
rect 431206 222618 437546 222854
rect 438102 222938 461690 223174
rect 461926 222938 473546 223174
rect 438102 222854 473546 222938
rect 438102 222618 461690 222854
rect 461926 222618 473546 222854
rect 474102 222938 492410 223174
rect 492646 222938 509546 223174
rect 474102 222854 509546 222938
rect 474102 222618 492410 222854
rect 492646 222618 509546 222854
rect 510102 222938 523130 223174
rect 523366 222938 545546 223174
rect 510102 222854 545546 222938
rect 510102 222618 523130 222854
rect 523366 222618 545546 222854
rect 546102 222938 553850 223174
rect 554086 222938 581546 223174
rect 546102 222854 581546 222938
rect 546102 222618 553850 222854
rect 554086 222618 581546 222854
rect 582102 222618 586302 223174
rect 586858 222618 592650 223174
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 218898 -1974 219454
rect -1418 218898 1826 219454
rect 2382 219218 16250 219454
rect 16486 219218 37826 219454
rect 2382 219134 37826 219218
rect 2382 218898 16250 219134
rect 16486 218898 37826 219134
rect 38382 219218 46970 219454
rect 47206 219218 73826 219454
rect 38382 219134 73826 219218
rect 38382 218898 46970 219134
rect 47206 218898 73826 219134
rect 74382 219218 77690 219454
rect 77926 219218 108410 219454
rect 108646 219218 109826 219454
rect 74382 219134 109826 219218
rect 74382 218898 77690 219134
rect 77926 218898 108410 219134
rect 108646 218898 109826 219134
rect 110382 219218 139130 219454
rect 139366 219218 145826 219454
rect 110382 219134 145826 219218
rect 110382 218898 139130 219134
rect 139366 218898 145826 219134
rect 146382 219218 169850 219454
rect 170086 219218 181826 219454
rect 146382 219134 181826 219218
rect 146382 218898 169850 219134
rect 170086 218898 181826 219134
rect 182382 219218 200570 219454
rect 200806 219218 217826 219454
rect 182382 219134 217826 219218
rect 182382 218898 200570 219134
rect 200806 218898 217826 219134
rect 218382 219218 231290 219454
rect 231526 219218 253826 219454
rect 218382 219134 253826 219218
rect 218382 218898 231290 219134
rect 231526 218898 253826 219134
rect 254382 219218 262010 219454
rect 262246 219218 289826 219454
rect 254382 219134 289826 219218
rect 254382 218898 262010 219134
rect 262246 218898 289826 219134
rect 290382 219218 292730 219454
rect 292966 219218 323450 219454
rect 323686 219218 325826 219454
rect 290382 219134 325826 219218
rect 290382 218898 292730 219134
rect 292966 218898 323450 219134
rect 323686 218898 325826 219134
rect 326382 219218 354170 219454
rect 354406 219218 361826 219454
rect 326382 219134 361826 219218
rect 326382 218898 354170 219134
rect 354406 218898 361826 219134
rect 362382 219218 384890 219454
rect 385126 219218 397826 219454
rect 362382 219134 397826 219218
rect 362382 218898 384890 219134
rect 385126 218898 397826 219134
rect 398382 219218 415610 219454
rect 415846 219218 433826 219454
rect 398382 219134 433826 219218
rect 398382 218898 415610 219134
rect 415846 218898 433826 219134
rect 434382 219218 446330 219454
rect 446566 219218 469826 219454
rect 434382 219134 469826 219218
rect 434382 218898 446330 219134
rect 446566 218898 469826 219134
rect 470382 219218 477050 219454
rect 477286 219218 505826 219454
rect 470382 219134 505826 219218
rect 470382 218898 477050 219134
rect 477286 218898 505826 219134
rect 506382 219218 507770 219454
rect 508006 219218 538490 219454
rect 538726 219218 541826 219454
rect 506382 219134 541826 219218
rect 506382 218898 507770 219134
rect 508006 218898 538490 219134
rect 538726 218898 541826 219134
rect 542382 219218 569210 219454
rect 569446 219218 577826 219454
rect 542382 219134 577826 219218
rect 542382 218898 569210 219134
rect 569446 218898 577826 219134
rect 578382 218898 585342 219454
rect 585898 218898 592650 219454
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 208938 -8694 209494
rect -8138 208938 27866 209494
rect 28422 208938 63866 209494
rect 64422 208938 99866 209494
rect 100422 208938 135866 209494
rect 136422 208938 171866 209494
rect 172422 208938 207866 209494
rect 208422 208938 243866 209494
rect 244422 208938 279866 209494
rect 280422 208938 315866 209494
rect 316422 208938 351866 209494
rect 352422 208938 387866 209494
rect 388422 208938 423866 209494
rect 424422 208938 459866 209494
rect 460422 208938 495866 209494
rect 496422 208938 531866 209494
rect 532422 208938 567866 209494
rect 568422 208938 592062 209494
rect 592618 208938 592650 209494
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205218 -7734 205774
rect -7178 205218 24146 205774
rect 24702 205218 60146 205774
rect 60702 205218 96146 205774
rect 96702 205218 132146 205774
rect 132702 205218 168146 205774
rect 168702 205218 204146 205774
rect 204702 205218 240146 205774
rect 240702 205218 276146 205774
rect 276702 205218 312146 205774
rect 312702 205218 348146 205774
rect 348702 205218 420146 205774
rect 420702 205218 456146 205774
rect 456702 205218 528146 205774
rect 528702 205218 564146 205774
rect 564702 205218 591102 205774
rect 591658 205218 592650 205774
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201498 -6774 202054
rect -6218 201498 20426 202054
rect 20982 201498 56426 202054
rect 56982 201498 128426 202054
rect 128982 201498 164426 202054
rect 164982 201498 236426 202054
rect 236982 201498 272426 202054
rect 272982 201498 344426 202054
rect 344982 201498 380426 202054
rect 380982 201498 416426 202054
rect 416982 201498 452426 202054
rect 452982 201498 488426 202054
rect 488982 201498 524426 202054
rect 524982 201498 560426 202054
rect 560982 201498 590142 202054
rect 590698 201498 592650 202054
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 197778 -5814 198334
rect -5258 197778 16706 198334
rect 17262 197778 52706 198334
rect 53262 197778 88706 198334
rect 89262 197778 124706 198334
rect 125262 197778 160706 198334
rect 161262 197778 196706 198334
rect 197262 197778 232706 198334
rect 233262 197778 268706 198334
rect 269262 197778 304706 198334
rect 305262 197778 340706 198334
rect 341262 197778 376706 198334
rect 377262 197778 412706 198334
rect 413262 197778 448706 198334
rect 449262 197778 484706 198334
rect 485262 197778 520706 198334
rect 521262 197778 556706 198334
rect 557262 197778 589182 198334
rect 589738 197778 592650 198334
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194058 -4854 194614
rect -4298 194058 12986 194614
rect 13542 194058 48986 194614
rect 49542 194058 84986 194614
rect 85542 194058 120986 194614
rect 121542 194058 156986 194614
rect 157542 194058 192986 194614
rect 193542 194058 228986 194614
rect 229542 194058 264986 194614
rect 265542 194058 300986 194614
rect 301542 194058 336986 194614
rect 337542 194058 372986 194614
rect 373542 194058 408986 194614
rect 409542 194058 444986 194614
rect 445542 194058 480986 194614
rect 481542 194058 516986 194614
rect 517542 194058 552986 194614
rect 553542 194058 588222 194614
rect 588778 194058 592650 194614
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190338 -3894 190894
rect -3338 190338 9266 190894
rect 9822 190338 45266 190894
rect 45822 190338 81266 190894
rect 81822 190338 117266 190894
rect 117822 190338 153266 190894
rect 153822 190338 189266 190894
rect 189822 190338 225266 190894
rect 225822 190338 297266 190894
rect 297822 190338 333266 190894
rect 333822 190338 405266 190894
rect 405822 190338 441266 190894
rect 441822 190338 513266 190894
rect 513822 190338 549266 190894
rect 549822 190338 587262 190894
rect 587818 190338 592650 190894
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186618 -2934 187174
rect -2378 186618 5546 187174
rect 6102 186938 31610 187174
rect 31846 186938 41546 187174
rect 6102 186854 41546 186938
rect 6102 186618 31610 186854
rect 31846 186618 41546 186854
rect 42102 186938 62330 187174
rect 62566 186938 93050 187174
rect 93286 186938 113546 187174
rect 42102 186854 113546 186938
rect 42102 186618 62330 186854
rect 62566 186618 93050 186854
rect 93286 186618 113546 186854
rect 114102 186938 123770 187174
rect 124006 186938 149546 187174
rect 114102 186854 149546 186938
rect 114102 186618 123770 186854
rect 124006 186618 149546 186854
rect 150102 186938 154490 187174
rect 154726 186938 185210 187174
rect 185446 186938 215930 187174
rect 216166 186938 221546 187174
rect 150102 186854 221546 186938
rect 150102 186618 154490 186854
rect 154726 186618 185210 186854
rect 185446 186618 215930 186854
rect 216166 186618 221546 186854
rect 222102 186938 246650 187174
rect 246886 186938 257546 187174
rect 222102 186854 257546 186938
rect 222102 186618 246650 186854
rect 246886 186618 257546 186854
rect 258102 186938 277370 187174
rect 277606 186938 293546 187174
rect 258102 186854 293546 186938
rect 258102 186618 277370 186854
rect 277606 186618 293546 186854
rect 294102 186938 308090 187174
rect 308326 186938 329546 187174
rect 294102 186854 329546 186938
rect 294102 186618 308090 186854
rect 308326 186618 329546 186854
rect 330102 186938 338810 187174
rect 339046 186938 365546 187174
rect 330102 186854 365546 186938
rect 330102 186618 338810 186854
rect 339046 186618 365546 186854
rect 366102 186938 369530 187174
rect 369766 186938 400250 187174
rect 400486 186938 401546 187174
rect 366102 186854 401546 186938
rect 366102 186618 369530 186854
rect 369766 186618 400250 186854
rect 400486 186618 401546 186854
rect 402102 186938 430970 187174
rect 431206 186938 437546 187174
rect 402102 186854 437546 186938
rect 402102 186618 430970 186854
rect 431206 186618 437546 186854
rect 438102 186938 461690 187174
rect 461926 186938 473546 187174
rect 438102 186854 473546 186938
rect 438102 186618 461690 186854
rect 461926 186618 473546 186854
rect 474102 186938 492410 187174
rect 492646 186938 509546 187174
rect 474102 186854 509546 186938
rect 474102 186618 492410 186854
rect 492646 186618 509546 186854
rect 510102 186938 523130 187174
rect 523366 186938 545546 187174
rect 510102 186854 545546 186938
rect 510102 186618 523130 186854
rect 523366 186618 545546 186854
rect 546102 186938 553850 187174
rect 554086 186938 581546 187174
rect 546102 186854 581546 186938
rect 546102 186618 553850 186854
rect 554086 186618 581546 186854
rect 582102 186618 586302 187174
rect 586858 186618 592650 187174
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 182898 -1974 183454
rect -1418 182898 1826 183454
rect 2382 183218 16250 183454
rect 16486 183218 37826 183454
rect 2382 183134 37826 183218
rect 2382 182898 16250 183134
rect 16486 182898 37826 183134
rect 38382 183218 46970 183454
rect 47206 183218 73826 183454
rect 38382 183134 73826 183218
rect 38382 182898 46970 183134
rect 47206 182898 73826 183134
rect 74382 183218 77690 183454
rect 77926 183218 108410 183454
rect 108646 183218 109826 183454
rect 74382 183134 109826 183218
rect 74382 182898 77690 183134
rect 77926 182898 108410 183134
rect 108646 182898 109826 183134
rect 110382 183218 139130 183454
rect 139366 183218 145826 183454
rect 110382 183134 145826 183218
rect 110382 182898 139130 183134
rect 139366 182898 145826 183134
rect 146382 183218 169850 183454
rect 170086 183218 181826 183454
rect 146382 183134 181826 183218
rect 146382 182898 169850 183134
rect 170086 182898 181826 183134
rect 182382 183218 200570 183454
rect 200806 183218 217826 183454
rect 182382 183134 217826 183218
rect 182382 182898 200570 183134
rect 200806 182898 217826 183134
rect 218382 183218 231290 183454
rect 231526 183218 253826 183454
rect 218382 183134 253826 183218
rect 218382 182898 231290 183134
rect 231526 182898 253826 183134
rect 254382 183218 262010 183454
rect 262246 183218 289826 183454
rect 254382 183134 289826 183218
rect 254382 182898 262010 183134
rect 262246 182898 289826 183134
rect 290382 183218 292730 183454
rect 292966 183218 323450 183454
rect 323686 183218 325826 183454
rect 290382 183134 325826 183218
rect 290382 182898 292730 183134
rect 292966 182898 323450 183134
rect 323686 182898 325826 183134
rect 326382 183218 354170 183454
rect 354406 183218 361826 183454
rect 326382 183134 361826 183218
rect 326382 182898 354170 183134
rect 354406 182898 361826 183134
rect 362382 183218 384890 183454
rect 385126 183218 397826 183454
rect 362382 183134 397826 183218
rect 362382 182898 384890 183134
rect 385126 182898 397826 183134
rect 398382 183218 415610 183454
rect 415846 183218 433826 183454
rect 398382 183134 433826 183218
rect 398382 182898 415610 183134
rect 415846 182898 433826 183134
rect 434382 183218 446330 183454
rect 446566 183218 469826 183454
rect 434382 183134 469826 183218
rect 434382 182898 446330 183134
rect 446566 182898 469826 183134
rect 470382 183218 477050 183454
rect 477286 183218 505826 183454
rect 470382 183134 505826 183218
rect 470382 182898 477050 183134
rect 477286 182898 505826 183134
rect 506382 183218 507770 183454
rect 508006 183218 538490 183454
rect 538726 183218 541826 183454
rect 506382 183134 541826 183218
rect 506382 182898 507770 183134
rect 508006 182898 538490 183134
rect 538726 182898 541826 183134
rect 542382 183218 569210 183454
rect 569446 183218 577826 183454
rect 542382 183134 577826 183218
rect 542382 182898 569210 183134
rect 569446 182898 577826 183134
rect 578382 182898 585342 183454
rect 585898 182898 592650 183454
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 172938 -8694 173494
rect -8138 172938 27866 173494
rect 28422 172938 63866 173494
rect 64422 172938 99866 173494
rect 100422 172938 135866 173494
rect 136422 172938 171866 173494
rect 172422 172938 207866 173494
rect 208422 172938 243866 173494
rect 244422 172938 279866 173494
rect 280422 172938 315866 173494
rect 316422 172938 351866 173494
rect 352422 172938 387866 173494
rect 388422 172938 423866 173494
rect 424422 172938 459866 173494
rect 460422 172938 495866 173494
rect 496422 172938 531866 173494
rect 532422 172938 567866 173494
rect 568422 172938 592062 173494
rect 592618 172938 592650 173494
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169218 -7734 169774
rect -7178 169218 24146 169774
rect 24702 169218 60146 169774
rect 60702 169218 96146 169774
rect 96702 169218 132146 169774
rect 132702 169218 168146 169774
rect 168702 169218 204146 169774
rect 204702 169218 240146 169774
rect 240702 169218 276146 169774
rect 276702 169218 312146 169774
rect 312702 169218 348146 169774
rect 348702 169218 420146 169774
rect 420702 169218 456146 169774
rect 456702 169218 528146 169774
rect 528702 169218 564146 169774
rect 564702 169218 591102 169774
rect 591658 169218 592650 169774
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165498 -6774 166054
rect -6218 165498 20426 166054
rect 20982 165498 56426 166054
rect 56982 165498 128426 166054
rect 128982 165498 164426 166054
rect 164982 165498 236426 166054
rect 236982 165498 272426 166054
rect 272982 165498 344426 166054
rect 344982 165498 380426 166054
rect 380982 165498 416426 166054
rect 416982 165498 452426 166054
rect 452982 165498 488426 166054
rect 488982 165498 524426 166054
rect 524982 165498 560426 166054
rect 560982 165498 590142 166054
rect 590698 165498 592650 166054
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 161778 -5814 162334
rect -5258 161778 16706 162334
rect 17262 161778 52706 162334
rect 53262 161778 88706 162334
rect 89262 161778 124706 162334
rect 125262 161778 160706 162334
rect 161262 161778 196706 162334
rect 197262 161778 232706 162334
rect 233262 161778 268706 162334
rect 269262 161778 304706 162334
rect 305262 161778 340706 162334
rect 341262 161778 376706 162334
rect 377262 161778 412706 162334
rect 413262 161778 448706 162334
rect 449262 161778 484706 162334
rect 485262 161778 520706 162334
rect 521262 161778 556706 162334
rect 557262 161778 589182 162334
rect 589738 161778 592650 162334
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158058 -4854 158614
rect -4298 158058 12986 158614
rect 13542 158058 48986 158614
rect 49542 158058 84986 158614
rect 85542 158058 120986 158614
rect 121542 158058 156986 158614
rect 157542 158058 192986 158614
rect 193542 158058 228986 158614
rect 229542 158058 264986 158614
rect 265542 158058 300986 158614
rect 301542 158058 336986 158614
rect 337542 158058 372986 158614
rect 373542 158058 408986 158614
rect 409542 158058 444986 158614
rect 445542 158058 480986 158614
rect 481542 158058 516986 158614
rect 517542 158058 552986 158614
rect 553542 158058 588222 158614
rect 588778 158058 592650 158614
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154338 -3894 154894
rect -3338 154338 9266 154894
rect 9822 154338 45266 154894
rect 45822 154338 81266 154894
rect 81822 154338 117266 154894
rect 117822 154338 153266 154894
rect 153822 154338 189266 154894
rect 189822 154338 225266 154894
rect 225822 154338 297266 154894
rect 297822 154338 333266 154894
rect 333822 154338 405266 154894
rect 405822 154338 441266 154894
rect 441822 154338 513266 154894
rect 513822 154338 549266 154894
rect 549822 154338 587262 154894
rect 587818 154338 592650 154894
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150618 -2934 151174
rect -2378 150618 5546 151174
rect 6102 150938 31610 151174
rect 31846 150938 41546 151174
rect 6102 150854 41546 150938
rect 6102 150618 31610 150854
rect 31846 150618 41546 150854
rect 42102 150938 62330 151174
rect 62566 150938 93050 151174
rect 93286 150938 113546 151174
rect 42102 150854 113546 150938
rect 42102 150618 62330 150854
rect 62566 150618 93050 150854
rect 93286 150618 113546 150854
rect 114102 150938 123770 151174
rect 124006 150938 149546 151174
rect 114102 150854 149546 150938
rect 114102 150618 123770 150854
rect 124006 150618 149546 150854
rect 150102 150938 154490 151174
rect 154726 150938 185210 151174
rect 185446 150938 215930 151174
rect 216166 150938 221546 151174
rect 150102 150854 221546 150938
rect 150102 150618 154490 150854
rect 154726 150618 185210 150854
rect 185446 150618 215930 150854
rect 216166 150618 221546 150854
rect 222102 150938 246650 151174
rect 246886 150938 257546 151174
rect 222102 150854 257546 150938
rect 222102 150618 246650 150854
rect 246886 150618 257546 150854
rect 258102 150938 277370 151174
rect 277606 150938 293546 151174
rect 258102 150854 293546 150938
rect 258102 150618 277370 150854
rect 277606 150618 293546 150854
rect 294102 150938 308090 151174
rect 308326 150938 329546 151174
rect 294102 150854 329546 150938
rect 294102 150618 308090 150854
rect 308326 150618 329546 150854
rect 330102 150938 338810 151174
rect 339046 150938 365546 151174
rect 330102 150854 365546 150938
rect 330102 150618 338810 150854
rect 339046 150618 365546 150854
rect 366102 150938 369530 151174
rect 369766 150938 400250 151174
rect 400486 150938 401546 151174
rect 366102 150854 401546 150938
rect 366102 150618 369530 150854
rect 369766 150618 400250 150854
rect 400486 150618 401546 150854
rect 402102 150938 430970 151174
rect 431206 150938 437546 151174
rect 402102 150854 437546 150938
rect 402102 150618 430970 150854
rect 431206 150618 437546 150854
rect 438102 150938 461690 151174
rect 461926 150938 473546 151174
rect 438102 150854 473546 150938
rect 438102 150618 461690 150854
rect 461926 150618 473546 150854
rect 474102 150938 492410 151174
rect 492646 150938 509546 151174
rect 474102 150854 509546 150938
rect 474102 150618 492410 150854
rect 492646 150618 509546 150854
rect 510102 150938 523130 151174
rect 523366 150938 545546 151174
rect 510102 150854 545546 150938
rect 510102 150618 523130 150854
rect 523366 150618 545546 150854
rect 546102 150938 553850 151174
rect 554086 150938 581546 151174
rect 546102 150854 581546 150938
rect 546102 150618 553850 150854
rect 554086 150618 581546 150854
rect 582102 150618 586302 151174
rect 586858 150618 592650 151174
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 146898 -1974 147454
rect -1418 146898 1826 147454
rect 2382 147218 16250 147454
rect 16486 147218 37826 147454
rect 2382 147134 37826 147218
rect 2382 146898 16250 147134
rect 16486 146898 37826 147134
rect 38382 147218 46970 147454
rect 47206 147218 73826 147454
rect 38382 147134 73826 147218
rect 38382 146898 46970 147134
rect 47206 146898 73826 147134
rect 74382 147218 77690 147454
rect 77926 147218 108410 147454
rect 108646 147218 109826 147454
rect 74382 147134 109826 147218
rect 74382 146898 77690 147134
rect 77926 146898 108410 147134
rect 108646 146898 109826 147134
rect 110382 147218 139130 147454
rect 139366 147218 145826 147454
rect 110382 147134 145826 147218
rect 110382 146898 139130 147134
rect 139366 146898 145826 147134
rect 146382 147218 169850 147454
rect 170086 147218 181826 147454
rect 146382 147134 181826 147218
rect 146382 146898 169850 147134
rect 170086 146898 181826 147134
rect 182382 147218 200570 147454
rect 200806 147218 217826 147454
rect 182382 147134 217826 147218
rect 182382 146898 200570 147134
rect 200806 146898 217826 147134
rect 218382 147218 231290 147454
rect 231526 147218 253826 147454
rect 218382 147134 253826 147218
rect 218382 146898 231290 147134
rect 231526 146898 253826 147134
rect 254382 147218 262010 147454
rect 262246 147218 289826 147454
rect 254382 147134 289826 147218
rect 254382 146898 262010 147134
rect 262246 146898 289826 147134
rect 290382 147218 292730 147454
rect 292966 147218 323450 147454
rect 323686 147218 325826 147454
rect 290382 147134 325826 147218
rect 290382 146898 292730 147134
rect 292966 146898 323450 147134
rect 323686 146898 325826 147134
rect 326382 147218 354170 147454
rect 354406 147218 361826 147454
rect 326382 147134 361826 147218
rect 326382 146898 354170 147134
rect 354406 146898 361826 147134
rect 362382 147218 384890 147454
rect 385126 147218 397826 147454
rect 362382 147134 397826 147218
rect 362382 146898 384890 147134
rect 385126 146898 397826 147134
rect 398382 147218 415610 147454
rect 415846 147218 433826 147454
rect 398382 147134 433826 147218
rect 398382 146898 415610 147134
rect 415846 146898 433826 147134
rect 434382 147218 446330 147454
rect 446566 147218 469826 147454
rect 434382 147134 469826 147218
rect 434382 146898 446330 147134
rect 446566 146898 469826 147134
rect 470382 147218 477050 147454
rect 477286 147218 505826 147454
rect 470382 147134 505826 147218
rect 470382 146898 477050 147134
rect 477286 146898 505826 147134
rect 506382 147218 507770 147454
rect 508006 147218 538490 147454
rect 538726 147218 541826 147454
rect 506382 147134 541826 147218
rect 506382 146898 507770 147134
rect 508006 146898 538490 147134
rect 538726 146898 541826 147134
rect 542382 147218 569210 147454
rect 569446 147218 577826 147454
rect 542382 147134 577826 147218
rect 542382 146898 569210 147134
rect 569446 146898 577826 147134
rect 578382 146898 585342 147454
rect 585898 146898 592650 147454
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 136938 -8694 137494
rect -8138 136938 27866 137494
rect 28422 136938 63866 137494
rect 64422 136938 99866 137494
rect 100422 136938 135866 137494
rect 136422 136938 171866 137494
rect 172422 136938 207866 137494
rect 208422 136938 243866 137494
rect 244422 136938 279866 137494
rect 280422 136938 315866 137494
rect 316422 136938 351866 137494
rect 352422 136938 387866 137494
rect 388422 136938 423866 137494
rect 424422 136938 459866 137494
rect 460422 136938 495866 137494
rect 496422 136938 531866 137494
rect 532422 136938 567866 137494
rect 568422 136938 592062 137494
rect 592618 136938 592650 137494
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133218 -7734 133774
rect -7178 133218 24146 133774
rect 24702 133218 60146 133774
rect 60702 133218 96146 133774
rect 96702 133218 132146 133774
rect 132702 133218 168146 133774
rect 168702 133218 204146 133774
rect 204702 133218 240146 133774
rect 240702 133218 276146 133774
rect 276702 133218 312146 133774
rect 312702 133218 348146 133774
rect 348702 133218 420146 133774
rect 420702 133218 456146 133774
rect 456702 133218 528146 133774
rect 528702 133218 564146 133774
rect 564702 133218 591102 133774
rect 591658 133218 592650 133774
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129498 -6774 130054
rect -6218 129498 20426 130054
rect 20982 129498 56426 130054
rect 56982 129498 128426 130054
rect 128982 129498 164426 130054
rect 164982 129498 236426 130054
rect 236982 129498 272426 130054
rect 272982 129498 344426 130054
rect 344982 129498 380426 130054
rect 380982 129498 416426 130054
rect 416982 129498 452426 130054
rect 452982 129498 488426 130054
rect 488982 129498 524426 130054
rect 524982 129498 560426 130054
rect 560982 129498 590142 130054
rect 590698 129498 592650 130054
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 125778 -5814 126334
rect -5258 125778 16706 126334
rect 17262 125778 52706 126334
rect 53262 125778 88706 126334
rect 89262 125778 124706 126334
rect 125262 125778 160706 126334
rect 161262 125778 196706 126334
rect 197262 125778 232706 126334
rect 233262 125778 268706 126334
rect 269262 125778 304706 126334
rect 305262 125778 340706 126334
rect 341262 125778 376706 126334
rect 377262 125778 412706 126334
rect 413262 125778 448706 126334
rect 449262 125778 484706 126334
rect 485262 125778 520706 126334
rect 521262 125778 556706 126334
rect 557262 125778 589182 126334
rect 589738 125778 592650 126334
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122058 -4854 122614
rect -4298 122058 12986 122614
rect 13542 122058 48986 122614
rect 49542 122058 84986 122614
rect 85542 122058 120986 122614
rect 121542 122058 156986 122614
rect 157542 122058 192986 122614
rect 193542 122058 228986 122614
rect 229542 122058 264986 122614
rect 265542 122058 300986 122614
rect 301542 122058 336986 122614
rect 337542 122058 372986 122614
rect 373542 122058 408986 122614
rect 409542 122058 444986 122614
rect 445542 122058 480986 122614
rect 481542 122058 516986 122614
rect 517542 122058 552986 122614
rect 553542 122058 588222 122614
rect 588778 122058 592650 122614
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118338 -3894 118894
rect -3338 118338 9266 118894
rect 9822 118338 45266 118894
rect 45822 118338 81266 118894
rect 81822 118338 117266 118894
rect 117822 118338 153266 118894
rect 153822 118338 189266 118894
rect 189822 118338 225266 118894
rect 225822 118338 297266 118894
rect 297822 118338 333266 118894
rect 333822 118338 405266 118894
rect 405822 118338 441266 118894
rect 441822 118338 513266 118894
rect 513822 118338 549266 118894
rect 549822 118338 587262 118894
rect 587818 118338 592650 118894
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114618 -2934 115174
rect -2378 114618 5546 115174
rect 6102 114938 31610 115174
rect 31846 114938 41546 115174
rect 6102 114854 41546 114938
rect 6102 114618 31610 114854
rect 31846 114618 41546 114854
rect 42102 114938 62330 115174
rect 62566 114938 93050 115174
rect 93286 114938 113546 115174
rect 42102 114854 113546 114938
rect 42102 114618 62330 114854
rect 62566 114618 93050 114854
rect 93286 114618 113546 114854
rect 114102 114938 123770 115174
rect 124006 114938 149546 115174
rect 114102 114854 149546 114938
rect 114102 114618 123770 114854
rect 124006 114618 149546 114854
rect 150102 114938 154490 115174
rect 154726 114938 185210 115174
rect 185446 114938 215930 115174
rect 216166 114938 221546 115174
rect 150102 114854 221546 114938
rect 150102 114618 154490 114854
rect 154726 114618 185210 114854
rect 185446 114618 215930 114854
rect 216166 114618 221546 114854
rect 222102 114938 246650 115174
rect 246886 114938 257546 115174
rect 222102 114854 257546 114938
rect 222102 114618 246650 114854
rect 246886 114618 257546 114854
rect 258102 114938 277370 115174
rect 277606 114938 293546 115174
rect 258102 114854 293546 114938
rect 258102 114618 277370 114854
rect 277606 114618 293546 114854
rect 294102 114938 308090 115174
rect 308326 114938 329546 115174
rect 294102 114854 329546 114938
rect 294102 114618 308090 114854
rect 308326 114618 329546 114854
rect 330102 114938 338810 115174
rect 339046 114938 365546 115174
rect 330102 114854 365546 114938
rect 330102 114618 338810 114854
rect 339046 114618 365546 114854
rect 366102 114938 369530 115174
rect 369766 114938 400250 115174
rect 400486 114938 401546 115174
rect 366102 114854 401546 114938
rect 366102 114618 369530 114854
rect 369766 114618 400250 114854
rect 400486 114618 401546 114854
rect 402102 114938 430970 115174
rect 431206 114938 437546 115174
rect 402102 114854 437546 114938
rect 402102 114618 430970 114854
rect 431206 114618 437546 114854
rect 438102 114938 461690 115174
rect 461926 114938 473546 115174
rect 438102 114854 473546 114938
rect 438102 114618 461690 114854
rect 461926 114618 473546 114854
rect 474102 114938 492410 115174
rect 492646 114938 509546 115174
rect 474102 114854 509546 114938
rect 474102 114618 492410 114854
rect 492646 114618 509546 114854
rect 510102 114938 523130 115174
rect 523366 114938 545546 115174
rect 510102 114854 545546 114938
rect 510102 114618 523130 114854
rect 523366 114618 545546 114854
rect 546102 114938 553850 115174
rect 554086 114938 581546 115174
rect 546102 114854 581546 114938
rect 546102 114618 553850 114854
rect 554086 114618 581546 114854
rect 582102 114618 586302 115174
rect 586858 114618 592650 115174
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 110898 -1974 111454
rect -1418 110898 1826 111454
rect 2382 111218 16250 111454
rect 16486 111218 37826 111454
rect 2382 111134 37826 111218
rect 2382 110898 16250 111134
rect 16486 110898 37826 111134
rect 38382 111218 46970 111454
rect 47206 111218 73826 111454
rect 38382 111134 73826 111218
rect 38382 110898 46970 111134
rect 47206 110898 73826 111134
rect 74382 111218 77690 111454
rect 77926 111218 108410 111454
rect 108646 111218 109826 111454
rect 74382 111134 109826 111218
rect 74382 110898 77690 111134
rect 77926 110898 108410 111134
rect 108646 110898 109826 111134
rect 110382 111218 139130 111454
rect 139366 111218 145826 111454
rect 110382 111134 145826 111218
rect 110382 110898 139130 111134
rect 139366 110898 145826 111134
rect 146382 111218 169850 111454
rect 170086 111218 181826 111454
rect 146382 111134 181826 111218
rect 146382 110898 169850 111134
rect 170086 110898 181826 111134
rect 182382 111218 200570 111454
rect 200806 111218 217826 111454
rect 182382 111134 217826 111218
rect 182382 110898 200570 111134
rect 200806 110898 217826 111134
rect 218382 111218 231290 111454
rect 231526 111218 253826 111454
rect 218382 111134 253826 111218
rect 218382 110898 231290 111134
rect 231526 110898 253826 111134
rect 254382 111218 262010 111454
rect 262246 111218 289826 111454
rect 254382 111134 289826 111218
rect 254382 110898 262010 111134
rect 262246 110898 289826 111134
rect 290382 111218 292730 111454
rect 292966 111218 323450 111454
rect 323686 111218 325826 111454
rect 290382 111134 325826 111218
rect 290382 110898 292730 111134
rect 292966 110898 323450 111134
rect 323686 110898 325826 111134
rect 326382 111218 354170 111454
rect 354406 111218 361826 111454
rect 326382 111134 361826 111218
rect 326382 110898 354170 111134
rect 354406 110898 361826 111134
rect 362382 111218 384890 111454
rect 385126 111218 397826 111454
rect 362382 111134 397826 111218
rect 362382 110898 384890 111134
rect 385126 110898 397826 111134
rect 398382 111218 415610 111454
rect 415846 111218 433826 111454
rect 398382 111134 433826 111218
rect 398382 110898 415610 111134
rect 415846 110898 433826 111134
rect 434382 111218 446330 111454
rect 446566 111218 469826 111454
rect 434382 111134 469826 111218
rect 434382 110898 446330 111134
rect 446566 110898 469826 111134
rect 470382 111218 477050 111454
rect 477286 111218 505826 111454
rect 470382 111134 505826 111218
rect 470382 110898 477050 111134
rect 477286 110898 505826 111134
rect 506382 111218 507770 111454
rect 508006 111218 538490 111454
rect 538726 111218 541826 111454
rect 506382 111134 541826 111218
rect 506382 110898 507770 111134
rect 508006 110898 538490 111134
rect 538726 110898 541826 111134
rect 542382 111218 569210 111454
rect 569446 111218 577826 111454
rect 542382 111134 577826 111218
rect 542382 110898 569210 111134
rect 569446 110898 577826 111134
rect 578382 110898 585342 111454
rect 585898 110898 592650 111454
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 100938 -8694 101494
rect -8138 100938 27866 101494
rect 28422 100938 63866 101494
rect 64422 100938 99866 101494
rect 100422 100938 135866 101494
rect 136422 100938 171866 101494
rect 172422 100938 207866 101494
rect 208422 100938 243866 101494
rect 244422 100938 279866 101494
rect 280422 100938 315866 101494
rect 316422 100938 351866 101494
rect 352422 100938 387866 101494
rect 388422 100938 423866 101494
rect 424422 100938 459866 101494
rect 460422 100938 495866 101494
rect 496422 100938 531866 101494
rect 532422 100938 567866 101494
rect 568422 100938 592062 101494
rect 592618 100938 592650 101494
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97218 -7734 97774
rect -7178 97218 24146 97774
rect 24702 97218 60146 97774
rect 60702 97218 96146 97774
rect 96702 97218 132146 97774
rect 132702 97218 168146 97774
rect 168702 97218 204146 97774
rect 204702 97218 240146 97774
rect 240702 97218 276146 97774
rect 276702 97218 312146 97774
rect 312702 97218 348146 97774
rect 348702 97218 420146 97774
rect 420702 97218 456146 97774
rect 456702 97218 528146 97774
rect 528702 97218 564146 97774
rect 564702 97218 591102 97774
rect 591658 97218 592650 97774
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93498 -6774 94054
rect -6218 93498 20426 94054
rect 20982 93498 56426 94054
rect 56982 93498 128426 94054
rect 128982 93498 164426 94054
rect 164982 93498 236426 94054
rect 236982 93498 272426 94054
rect 272982 93498 344426 94054
rect 344982 93498 380426 94054
rect 380982 93498 416426 94054
rect 416982 93498 452426 94054
rect 452982 93498 488426 94054
rect 488982 93498 524426 94054
rect 524982 93498 560426 94054
rect 560982 93498 590142 94054
rect 590698 93498 592650 94054
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 89778 -5814 90334
rect -5258 89778 16706 90334
rect 17262 89778 52706 90334
rect 53262 89778 88706 90334
rect 89262 89778 124706 90334
rect 125262 89778 160706 90334
rect 161262 89778 196706 90334
rect 197262 89778 232706 90334
rect 233262 89778 268706 90334
rect 269262 89778 304706 90334
rect 305262 89778 340706 90334
rect 341262 89778 376706 90334
rect 377262 89778 412706 90334
rect 413262 89778 448706 90334
rect 449262 89778 484706 90334
rect 485262 89778 520706 90334
rect 521262 89778 556706 90334
rect 557262 89778 589182 90334
rect 589738 89778 592650 90334
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86058 -4854 86614
rect -4298 86058 12986 86614
rect 13542 86058 48986 86614
rect 49542 86058 84986 86614
rect 85542 86058 120986 86614
rect 121542 86058 156986 86614
rect 157542 86058 192986 86614
rect 193542 86058 228986 86614
rect 229542 86058 264986 86614
rect 265542 86058 300986 86614
rect 301542 86058 336986 86614
rect 337542 86058 372986 86614
rect 373542 86058 408986 86614
rect 409542 86058 444986 86614
rect 445542 86058 480986 86614
rect 481542 86058 516986 86614
rect 517542 86058 552986 86614
rect 553542 86058 588222 86614
rect 588778 86058 592650 86614
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82338 -3894 82894
rect -3338 82338 9266 82894
rect 9822 82338 45266 82894
rect 45822 82338 81266 82894
rect 81822 82338 117266 82894
rect 117822 82338 153266 82894
rect 153822 82338 189266 82894
rect 189822 82338 225266 82894
rect 225822 82338 297266 82894
rect 297822 82338 333266 82894
rect 333822 82338 405266 82894
rect 405822 82338 441266 82894
rect 441822 82338 513266 82894
rect 513822 82338 549266 82894
rect 549822 82338 587262 82894
rect 587818 82338 592650 82894
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78618 -2934 79174
rect -2378 78618 5546 79174
rect 6102 78938 31610 79174
rect 31846 78938 41546 79174
rect 6102 78854 41546 78938
rect 6102 78618 31610 78854
rect 31846 78618 41546 78854
rect 42102 78938 62330 79174
rect 62566 78938 93050 79174
rect 93286 78938 113546 79174
rect 42102 78854 113546 78938
rect 42102 78618 62330 78854
rect 62566 78618 93050 78854
rect 93286 78618 113546 78854
rect 114102 78938 123770 79174
rect 124006 78938 149546 79174
rect 114102 78854 149546 78938
rect 114102 78618 123770 78854
rect 124006 78618 149546 78854
rect 150102 78938 154490 79174
rect 154726 78938 185210 79174
rect 185446 78938 215930 79174
rect 216166 78938 221546 79174
rect 150102 78854 221546 78938
rect 150102 78618 154490 78854
rect 154726 78618 185210 78854
rect 185446 78618 215930 78854
rect 216166 78618 221546 78854
rect 222102 78938 246650 79174
rect 246886 78938 257546 79174
rect 222102 78854 257546 78938
rect 222102 78618 246650 78854
rect 246886 78618 257546 78854
rect 258102 78938 277370 79174
rect 277606 78938 293546 79174
rect 258102 78854 293546 78938
rect 258102 78618 277370 78854
rect 277606 78618 293546 78854
rect 294102 78938 308090 79174
rect 308326 78938 329546 79174
rect 294102 78854 329546 78938
rect 294102 78618 308090 78854
rect 308326 78618 329546 78854
rect 330102 78938 338810 79174
rect 339046 78938 365546 79174
rect 330102 78854 365546 78938
rect 330102 78618 338810 78854
rect 339046 78618 365546 78854
rect 366102 78938 369530 79174
rect 369766 78938 400250 79174
rect 400486 78938 401546 79174
rect 366102 78854 401546 78938
rect 366102 78618 369530 78854
rect 369766 78618 400250 78854
rect 400486 78618 401546 78854
rect 402102 78938 430970 79174
rect 431206 78938 437546 79174
rect 402102 78854 437546 78938
rect 402102 78618 430970 78854
rect 431206 78618 437546 78854
rect 438102 78938 461690 79174
rect 461926 78938 473546 79174
rect 438102 78854 473546 78938
rect 438102 78618 461690 78854
rect 461926 78618 473546 78854
rect 474102 78938 492410 79174
rect 492646 78938 509546 79174
rect 474102 78854 509546 78938
rect 474102 78618 492410 78854
rect 492646 78618 509546 78854
rect 510102 78938 523130 79174
rect 523366 78938 545546 79174
rect 510102 78854 545546 78938
rect 510102 78618 523130 78854
rect 523366 78618 545546 78854
rect 546102 78938 553850 79174
rect 554086 78938 581546 79174
rect 546102 78854 581546 78938
rect 546102 78618 553850 78854
rect 554086 78618 581546 78854
rect 582102 78618 586302 79174
rect 586858 78618 592650 79174
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 74898 -1974 75454
rect -1418 74898 1826 75454
rect 2382 75218 16250 75454
rect 16486 75218 37826 75454
rect 2382 75134 37826 75218
rect 2382 74898 16250 75134
rect 16486 74898 37826 75134
rect 38382 75218 46970 75454
rect 47206 75218 73826 75454
rect 38382 75134 73826 75218
rect 38382 74898 46970 75134
rect 47206 74898 73826 75134
rect 74382 75218 77690 75454
rect 77926 75218 108410 75454
rect 108646 75218 109826 75454
rect 74382 75134 109826 75218
rect 74382 74898 77690 75134
rect 77926 74898 108410 75134
rect 108646 74898 109826 75134
rect 110382 75218 139130 75454
rect 139366 75218 145826 75454
rect 110382 75134 145826 75218
rect 110382 74898 139130 75134
rect 139366 74898 145826 75134
rect 146382 75218 169850 75454
rect 170086 75218 181826 75454
rect 146382 75134 181826 75218
rect 146382 74898 169850 75134
rect 170086 74898 181826 75134
rect 182382 75218 200570 75454
rect 200806 75218 217826 75454
rect 182382 75134 217826 75218
rect 182382 74898 200570 75134
rect 200806 74898 217826 75134
rect 218382 75218 231290 75454
rect 231526 75218 253826 75454
rect 218382 75134 253826 75218
rect 218382 74898 231290 75134
rect 231526 74898 253826 75134
rect 254382 75218 262010 75454
rect 262246 75218 289826 75454
rect 254382 75134 289826 75218
rect 254382 74898 262010 75134
rect 262246 74898 289826 75134
rect 290382 75218 292730 75454
rect 292966 75218 323450 75454
rect 323686 75218 325826 75454
rect 290382 75134 325826 75218
rect 290382 74898 292730 75134
rect 292966 74898 323450 75134
rect 323686 74898 325826 75134
rect 326382 75218 354170 75454
rect 354406 75218 361826 75454
rect 326382 75134 361826 75218
rect 326382 74898 354170 75134
rect 354406 74898 361826 75134
rect 362382 75218 384890 75454
rect 385126 75218 397826 75454
rect 362382 75134 397826 75218
rect 362382 74898 384890 75134
rect 385126 74898 397826 75134
rect 398382 75218 415610 75454
rect 415846 75218 433826 75454
rect 398382 75134 433826 75218
rect 398382 74898 415610 75134
rect 415846 74898 433826 75134
rect 434382 75218 446330 75454
rect 446566 75218 469826 75454
rect 434382 75134 469826 75218
rect 434382 74898 446330 75134
rect 446566 74898 469826 75134
rect 470382 75218 477050 75454
rect 477286 75218 505826 75454
rect 470382 75134 505826 75218
rect 470382 74898 477050 75134
rect 477286 74898 505826 75134
rect 506382 75218 507770 75454
rect 508006 75218 538490 75454
rect 538726 75218 541826 75454
rect 506382 75134 541826 75218
rect 506382 74898 507770 75134
rect 508006 74898 538490 75134
rect 538726 74898 541826 75134
rect 542382 75218 569210 75454
rect 569446 75218 577826 75454
rect 542382 75134 577826 75218
rect 542382 74898 569210 75134
rect 569446 74898 577826 75134
rect 578382 74898 585342 75454
rect 585898 74898 592650 75454
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 64938 -8694 65494
rect -8138 64938 27866 65494
rect 28422 64938 63866 65494
rect 64422 64938 99866 65494
rect 100422 64938 135866 65494
rect 136422 64938 171866 65494
rect 172422 64938 207866 65494
rect 208422 64938 243866 65494
rect 244422 64938 279866 65494
rect 280422 64938 315866 65494
rect 316422 64938 351866 65494
rect 352422 64938 387866 65494
rect 388422 64938 423866 65494
rect 424422 64938 459866 65494
rect 460422 64938 495866 65494
rect 496422 64938 531866 65494
rect 532422 64938 567866 65494
rect 568422 64938 592062 65494
rect 592618 64938 592650 65494
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61218 -7734 61774
rect -7178 61218 24146 61774
rect 24702 61218 60146 61774
rect 60702 61218 96146 61774
rect 96702 61218 132146 61774
rect 132702 61218 168146 61774
rect 168702 61218 204146 61774
rect 204702 61218 240146 61774
rect 240702 61218 276146 61774
rect 276702 61218 312146 61774
rect 312702 61218 348146 61774
rect 348702 61218 420146 61774
rect 420702 61218 456146 61774
rect 456702 61218 528146 61774
rect 528702 61218 564146 61774
rect 564702 61218 591102 61774
rect 591658 61218 592650 61774
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57498 -6774 58054
rect -6218 57498 20426 58054
rect 20982 57498 56426 58054
rect 56982 57498 128426 58054
rect 128982 57498 164426 58054
rect 164982 57498 236426 58054
rect 236982 57498 272426 58054
rect 272982 57498 344426 58054
rect 344982 57498 380426 58054
rect 380982 57498 416426 58054
rect 416982 57498 452426 58054
rect 452982 57498 488426 58054
rect 488982 57498 524426 58054
rect 524982 57498 560426 58054
rect 560982 57498 590142 58054
rect 590698 57498 592650 58054
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 53778 -5814 54334
rect -5258 53778 16706 54334
rect 17262 53778 52706 54334
rect 53262 53778 88706 54334
rect 89262 53778 124706 54334
rect 125262 53778 160706 54334
rect 161262 53778 196706 54334
rect 197262 53778 232706 54334
rect 233262 53778 268706 54334
rect 269262 53778 304706 54334
rect 305262 53778 340706 54334
rect 341262 53778 376706 54334
rect 377262 53778 412706 54334
rect 413262 53778 448706 54334
rect 449262 53778 484706 54334
rect 485262 53778 520706 54334
rect 521262 53778 556706 54334
rect 557262 53778 589182 54334
rect 589738 53778 592650 54334
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50058 -4854 50614
rect -4298 50058 12986 50614
rect 13542 50058 48986 50614
rect 49542 50058 84986 50614
rect 85542 50058 120986 50614
rect 121542 50058 156986 50614
rect 157542 50058 192986 50614
rect 193542 50058 228986 50614
rect 229542 50058 264986 50614
rect 265542 50058 300986 50614
rect 301542 50058 336986 50614
rect 337542 50058 372986 50614
rect 373542 50058 408986 50614
rect 409542 50058 444986 50614
rect 445542 50058 480986 50614
rect 481542 50058 516986 50614
rect 517542 50058 552986 50614
rect 553542 50058 588222 50614
rect 588778 50058 592650 50614
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46338 -3894 46894
rect -3338 46338 9266 46894
rect 9822 46338 45266 46894
rect 45822 46338 81266 46894
rect 81822 46338 117266 46894
rect 117822 46338 153266 46894
rect 153822 46338 189266 46894
rect 189822 46338 225266 46894
rect 225822 46338 297266 46894
rect 297822 46338 333266 46894
rect 333822 46338 405266 46894
rect 405822 46338 441266 46894
rect 441822 46338 513266 46894
rect 513822 46338 549266 46894
rect 549822 46338 587262 46894
rect 587818 46338 592650 46894
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42618 -2934 43174
rect -2378 42618 5546 43174
rect 6102 42938 31610 43174
rect 31846 42938 41546 43174
rect 6102 42854 41546 42938
rect 6102 42618 31610 42854
rect 31846 42618 41546 42854
rect 42102 42938 62330 43174
rect 62566 42938 93050 43174
rect 93286 42938 113546 43174
rect 42102 42854 113546 42938
rect 42102 42618 62330 42854
rect 62566 42618 93050 42854
rect 93286 42618 113546 42854
rect 114102 42938 123770 43174
rect 124006 42938 149546 43174
rect 114102 42854 149546 42938
rect 114102 42618 123770 42854
rect 124006 42618 149546 42854
rect 150102 42938 154490 43174
rect 154726 42938 185210 43174
rect 185446 42938 215930 43174
rect 216166 42938 221546 43174
rect 150102 42854 221546 42938
rect 150102 42618 154490 42854
rect 154726 42618 185210 42854
rect 185446 42618 215930 42854
rect 216166 42618 221546 42854
rect 222102 42938 246650 43174
rect 246886 42938 257546 43174
rect 222102 42854 257546 42938
rect 222102 42618 246650 42854
rect 246886 42618 257546 42854
rect 258102 42938 277370 43174
rect 277606 42938 293546 43174
rect 258102 42854 293546 42938
rect 258102 42618 277370 42854
rect 277606 42618 293546 42854
rect 294102 42938 308090 43174
rect 308326 42938 329546 43174
rect 294102 42854 329546 42938
rect 294102 42618 308090 42854
rect 308326 42618 329546 42854
rect 330102 42938 338810 43174
rect 339046 42938 365546 43174
rect 330102 42854 365546 42938
rect 330102 42618 338810 42854
rect 339046 42618 365546 42854
rect 366102 42938 369530 43174
rect 369766 42938 400250 43174
rect 400486 42938 401546 43174
rect 366102 42854 401546 42938
rect 366102 42618 369530 42854
rect 369766 42618 400250 42854
rect 400486 42618 401546 42854
rect 402102 42938 430970 43174
rect 431206 42938 437546 43174
rect 402102 42854 437546 42938
rect 402102 42618 430970 42854
rect 431206 42618 437546 42854
rect 438102 42938 461690 43174
rect 461926 42938 473546 43174
rect 438102 42854 473546 42938
rect 438102 42618 461690 42854
rect 461926 42618 473546 42854
rect 474102 42938 492410 43174
rect 492646 42938 509546 43174
rect 474102 42854 509546 42938
rect 474102 42618 492410 42854
rect 492646 42618 509546 42854
rect 510102 42938 523130 43174
rect 523366 42938 545546 43174
rect 510102 42854 545546 42938
rect 510102 42618 523130 42854
rect 523366 42618 545546 42854
rect 546102 42938 553850 43174
rect 554086 42938 581546 43174
rect 546102 42854 581546 42938
rect 546102 42618 553850 42854
rect 554086 42618 581546 42854
rect 582102 42618 586302 43174
rect 586858 42618 592650 43174
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 38898 -1974 39454
rect -1418 38898 1826 39454
rect 2382 39218 16250 39454
rect 16486 39218 37826 39454
rect 2382 39134 37826 39218
rect 2382 38898 16250 39134
rect 16486 38898 37826 39134
rect 38382 39218 46970 39454
rect 47206 39218 73826 39454
rect 38382 39134 73826 39218
rect 38382 38898 46970 39134
rect 47206 38898 73826 39134
rect 74382 39218 77690 39454
rect 77926 39218 108410 39454
rect 108646 39218 109826 39454
rect 74382 39134 109826 39218
rect 74382 38898 77690 39134
rect 77926 38898 108410 39134
rect 108646 38898 109826 39134
rect 110382 39218 139130 39454
rect 139366 39218 145826 39454
rect 110382 39134 145826 39218
rect 110382 38898 139130 39134
rect 139366 38898 145826 39134
rect 146382 39218 169850 39454
rect 170086 39218 181826 39454
rect 146382 39134 181826 39218
rect 146382 38898 169850 39134
rect 170086 38898 181826 39134
rect 182382 39218 200570 39454
rect 200806 39218 217826 39454
rect 182382 39134 217826 39218
rect 182382 38898 200570 39134
rect 200806 38898 217826 39134
rect 218382 39218 231290 39454
rect 231526 39218 253826 39454
rect 218382 39134 253826 39218
rect 218382 38898 231290 39134
rect 231526 38898 253826 39134
rect 254382 39218 262010 39454
rect 262246 39218 289826 39454
rect 254382 39134 289826 39218
rect 254382 38898 262010 39134
rect 262246 38898 289826 39134
rect 290382 39218 292730 39454
rect 292966 39218 323450 39454
rect 323686 39218 325826 39454
rect 290382 39134 325826 39218
rect 290382 38898 292730 39134
rect 292966 38898 323450 39134
rect 323686 38898 325826 39134
rect 326382 39218 354170 39454
rect 354406 39218 361826 39454
rect 326382 39134 361826 39218
rect 326382 38898 354170 39134
rect 354406 38898 361826 39134
rect 362382 39218 384890 39454
rect 385126 39218 397826 39454
rect 362382 39134 397826 39218
rect 362382 38898 384890 39134
rect 385126 38898 397826 39134
rect 398382 39218 415610 39454
rect 415846 39218 433826 39454
rect 398382 39134 433826 39218
rect 398382 38898 415610 39134
rect 415846 38898 433826 39134
rect 434382 39218 446330 39454
rect 446566 39218 469826 39454
rect 434382 39134 469826 39218
rect 434382 38898 446330 39134
rect 446566 38898 469826 39134
rect 470382 39218 477050 39454
rect 477286 39218 505826 39454
rect 470382 39134 505826 39218
rect 470382 38898 477050 39134
rect 477286 38898 505826 39134
rect 506382 39218 507770 39454
rect 508006 39218 538490 39454
rect 538726 39218 541826 39454
rect 506382 39134 541826 39218
rect 506382 38898 507770 39134
rect 508006 38898 538490 39134
rect 538726 38898 541826 39134
rect 542382 39218 569210 39454
rect 569446 39218 577826 39454
rect 542382 39134 577826 39218
rect 542382 38898 569210 39134
rect 569446 38898 577826 39134
rect 578382 38898 585342 39454
rect 585898 38898 592650 39454
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 28938 -8694 29494
rect -8138 28938 27866 29494
rect 28422 28938 63866 29494
rect 64422 28938 99866 29494
rect 100422 28938 135866 29494
rect 136422 28938 171866 29494
rect 172422 28938 207866 29494
rect 208422 28938 243866 29494
rect 244422 28938 279866 29494
rect 280422 28938 315866 29494
rect 316422 28938 351866 29494
rect 352422 28938 387866 29494
rect 388422 28938 423866 29494
rect 424422 28938 459866 29494
rect 460422 28938 495866 29494
rect 496422 28938 531866 29494
rect 532422 28938 567866 29494
rect 568422 28938 592062 29494
rect 592618 28938 592650 29494
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25218 -7734 25774
rect -7178 25218 24146 25774
rect 24702 25218 60146 25774
rect 60702 25218 96146 25774
rect 96702 25218 132146 25774
rect 132702 25218 168146 25774
rect 168702 25218 204146 25774
rect 204702 25218 240146 25774
rect 240702 25218 276146 25774
rect 276702 25218 312146 25774
rect 312702 25218 348146 25774
rect 348702 25218 420146 25774
rect 420702 25218 456146 25774
rect 456702 25218 528146 25774
rect 528702 25218 564146 25774
rect 564702 25218 591102 25774
rect 591658 25218 592650 25774
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21498 -6774 22054
rect -6218 21498 20426 22054
rect 20982 21498 56426 22054
rect 56982 21498 128426 22054
rect 128982 21498 164426 22054
rect 164982 21498 236426 22054
rect 236982 21498 272426 22054
rect 272982 21498 344426 22054
rect 344982 21498 380426 22054
rect 380982 21498 416426 22054
rect 416982 21498 452426 22054
rect 452982 21498 488426 22054
rect 488982 21498 524426 22054
rect 524982 21498 560426 22054
rect 560982 21498 590142 22054
rect 590698 21498 592650 22054
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 17778 -5814 18334
rect -5258 17778 16706 18334
rect 17262 17778 52706 18334
rect 53262 17778 88706 18334
rect 89262 17778 124706 18334
rect 125262 17778 160706 18334
rect 161262 17778 196706 18334
rect 197262 17778 232706 18334
rect 233262 17778 268706 18334
rect 269262 17778 304706 18334
rect 305262 17778 340706 18334
rect 341262 17778 376706 18334
rect 377262 17778 412706 18334
rect 413262 17778 448706 18334
rect 449262 17778 484706 18334
rect 485262 17778 520706 18334
rect 521262 17778 556706 18334
rect 557262 17778 589182 18334
rect 589738 17778 592650 18334
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14058 -4854 14614
rect -4298 14058 12986 14614
rect 13542 14058 48986 14614
rect 49542 14058 84986 14614
rect 85542 14058 120986 14614
rect 121542 14058 156986 14614
rect 157542 14058 192986 14614
rect 193542 14058 228986 14614
rect 229542 14058 264986 14614
rect 265542 14058 300986 14614
rect 301542 14058 336986 14614
rect 337542 14058 372986 14614
rect 373542 14058 408986 14614
rect 409542 14058 444986 14614
rect 445542 14058 480986 14614
rect 481542 14058 516986 14614
rect 517542 14058 552986 14614
rect 553542 14058 588222 14614
rect 588778 14058 592650 14614
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10338 -3894 10894
rect -3338 10338 9266 10894
rect 9822 10338 45266 10894
rect 45822 10338 81266 10894
rect 81822 10338 117266 10894
rect 117822 10338 153266 10894
rect 153822 10338 189266 10894
rect 189822 10338 225266 10894
rect 225822 10338 297266 10894
rect 297822 10338 333266 10894
rect 333822 10338 405266 10894
rect 405822 10338 441266 10894
rect 441822 10338 513266 10894
rect 513822 10338 549266 10894
rect 549822 10338 587262 10894
rect 587818 10338 592650 10894
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6618 -2934 7174
rect -2378 6618 5546 7174
rect 6102 6938 31610 7174
rect 31846 6938 41546 7174
rect 6102 6854 41546 6938
rect 6102 6618 31610 6854
rect 31846 6618 41546 6854
rect 42102 6938 62330 7174
rect 62566 6938 93050 7174
rect 93286 6938 113546 7174
rect 42102 6854 113546 6938
rect 42102 6618 62330 6854
rect 62566 6618 93050 6854
rect 93286 6618 113546 6854
rect 114102 6938 123770 7174
rect 124006 6938 149546 7174
rect 114102 6854 149546 6938
rect 114102 6618 123770 6854
rect 124006 6618 149546 6854
rect 150102 6938 154490 7174
rect 154726 6938 185210 7174
rect 185446 6938 215930 7174
rect 216166 6938 221546 7174
rect 150102 6854 221546 6938
rect 150102 6618 154490 6854
rect 154726 6618 185210 6854
rect 185446 6618 215930 6854
rect 216166 6618 221546 6854
rect 222102 6938 246650 7174
rect 246886 6938 257546 7174
rect 222102 6854 257546 6938
rect 222102 6618 246650 6854
rect 246886 6618 257546 6854
rect 258102 6938 277370 7174
rect 277606 6938 293546 7174
rect 258102 6854 293546 6938
rect 258102 6618 277370 6854
rect 277606 6618 293546 6854
rect 294102 6938 308090 7174
rect 308326 6938 329546 7174
rect 294102 6854 329546 6938
rect 294102 6618 308090 6854
rect 308326 6618 329546 6854
rect 330102 6938 338810 7174
rect 339046 6938 365546 7174
rect 330102 6854 365546 6938
rect 330102 6618 338810 6854
rect 339046 6618 365546 6854
rect 366102 6938 369530 7174
rect 369766 6938 400250 7174
rect 400486 6938 401546 7174
rect 366102 6854 401546 6938
rect 366102 6618 369530 6854
rect 369766 6618 400250 6854
rect 400486 6618 401546 6854
rect 402102 6938 430970 7174
rect 431206 6938 437546 7174
rect 402102 6854 437546 6938
rect 402102 6618 430970 6854
rect 431206 6618 437546 6854
rect 438102 6938 461690 7174
rect 461926 6938 473546 7174
rect 438102 6854 473546 6938
rect 438102 6618 461690 6854
rect 461926 6618 473546 6854
rect 474102 6938 492410 7174
rect 492646 6938 509546 7174
rect 474102 6854 509546 6938
rect 474102 6618 492410 6854
rect 492646 6618 509546 6854
rect 510102 6938 523130 7174
rect 523366 6938 545546 7174
rect 510102 6854 545546 6938
rect 510102 6618 523130 6854
rect 523366 6618 545546 6854
rect 546102 6938 553850 7174
rect 554086 6938 581546 7174
rect 546102 6854 581546 6938
rect 546102 6618 553850 6854
rect 554086 6618 581546 6854
rect 582102 6618 586302 7174
rect 586858 6618 592650 7174
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 2898 -1974 3454
rect -1418 2898 1826 3454
rect 2382 2898 37826 3454
rect 38382 2898 73826 3454
rect 74382 2898 109826 3454
rect 110382 2898 145826 3454
rect 146382 2898 181826 3454
rect 182382 2898 217826 3454
rect 218382 2898 253826 3454
rect 254382 2898 289826 3454
rect 290382 2898 325826 3454
rect 326382 2898 361826 3454
rect 362382 2898 397826 3454
rect 398382 2898 433826 3454
rect 434382 2898 469826 3454
rect 470382 2898 505826 3454
rect 506382 2898 541826 3454
rect 542382 2898 577826 3454
rect 578382 2898 585342 3454
rect 585898 2898 592650 3454
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -902 -1974 -346
rect -1418 -902 1826 -346
rect 2382 -902 37826 -346
rect 38382 -902 73826 -346
rect 74382 -902 109826 -346
rect 110382 -902 145826 -346
rect 146382 -902 181826 -346
rect 182382 -902 217826 -346
rect 218382 -902 253826 -346
rect 254382 -902 289826 -346
rect 290382 -902 325826 -346
rect 326382 -902 361826 -346
rect 362382 -902 397826 -346
rect 398382 -902 433826 -346
rect 434382 -902 469826 -346
rect 470382 -902 505826 -346
rect 506382 -902 541826 -346
rect 542382 -902 577826 -346
rect 578382 -902 585342 -346
rect 585898 -902 585930 -346
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1862 -2934 -1306
rect -2378 -1862 5546 -1306
rect 6102 -1862 41546 -1306
rect 42102 -1862 113546 -1306
rect 114102 -1862 149546 -1306
rect 150102 -1862 221546 -1306
rect 222102 -1862 257546 -1306
rect 258102 -1862 293546 -1306
rect 294102 -1862 329546 -1306
rect 330102 -1862 365546 -1306
rect 366102 -1862 401546 -1306
rect 402102 -1862 437546 -1306
rect 438102 -1862 473546 -1306
rect 474102 -1862 509546 -1306
rect 510102 -1862 545546 -1306
rect 546102 -1862 581546 -1306
rect 582102 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2822 -3894 -2266
rect -3338 -2822 9266 -2266
rect 9822 -2822 45266 -2266
rect 45822 -2822 81266 -2266
rect 81822 -2822 117266 -2266
rect 117822 -2822 153266 -2266
rect 153822 -2822 189266 -2266
rect 189822 -2822 225266 -2266
rect 225822 -2822 297266 -2266
rect 297822 -2822 333266 -2266
rect 333822 -2822 405266 -2266
rect 405822 -2822 441266 -2266
rect 441822 -2822 513266 -2266
rect 513822 -2822 549266 -2266
rect 549822 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3782 -4854 -3226
rect -4298 -3782 12986 -3226
rect 13542 -3782 48986 -3226
rect 49542 -3782 84986 -3226
rect 85542 -3782 120986 -3226
rect 121542 -3782 156986 -3226
rect 157542 -3782 192986 -3226
rect 193542 -3782 228986 -3226
rect 229542 -3782 264986 -3226
rect 265542 -3782 300986 -3226
rect 301542 -3782 336986 -3226
rect 337542 -3782 372986 -3226
rect 373542 -3782 408986 -3226
rect 409542 -3782 444986 -3226
rect 445542 -3782 480986 -3226
rect 481542 -3782 516986 -3226
rect 517542 -3782 552986 -3226
rect 553542 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4742 -5814 -4186
rect -5258 -4742 16706 -4186
rect 17262 -4742 52706 -4186
rect 53262 -4742 88706 -4186
rect 89262 -4742 124706 -4186
rect 125262 -4742 160706 -4186
rect 161262 -4742 196706 -4186
rect 197262 -4742 232706 -4186
rect 233262 -4742 268706 -4186
rect 269262 -4742 304706 -4186
rect 305262 -4742 340706 -4186
rect 341262 -4742 376706 -4186
rect 377262 -4742 412706 -4186
rect 413262 -4742 448706 -4186
rect 449262 -4742 484706 -4186
rect 485262 -4742 520706 -4186
rect 521262 -4742 556706 -4186
rect 557262 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5702 -6774 -5146
rect -6218 -5702 20426 -5146
rect 20982 -5702 56426 -5146
rect 56982 -5702 128426 -5146
rect 128982 -5702 164426 -5146
rect 164982 -5702 236426 -5146
rect 236982 -5702 272426 -5146
rect 272982 -5702 344426 -5146
rect 344982 -5702 380426 -5146
rect 380982 -5702 416426 -5146
rect 416982 -5702 452426 -5146
rect 452982 -5702 488426 -5146
rect 488982 -5702 524426 -5146
rect 524982 -5702 560426 -5146
rect 560982 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6662 -7734 -6106
rect -7178 -6662 24146 -6106
rect 24702 -6662 60146 -6106
rect 60702 -6662 96146 -6106
rect 96702 -6662 132146 -6106
rect 132702 -6662 168146 -6106
rect 168702 -6662 204146 -6106
rect 204702 -6662 240146 -6106
rect 240702 -6662 276146 -6106
rect 276702 -6662 312146 -6106
rect 312702 -6662 348146 -6106
rect 348702 -6662 420146 -6106
rect 420702 -6662 456146 -6106
rect 456702 -6662 528146 -6106
rect 528702 -6662 564146 -6106
rect 564702 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7622 -8694 -7066
rect -8138 -7622 27866 -7066
rect 28422 -7622 63866 -7066
rect 64422 -7622 99866 -7066
rect 100422 -7622 135866 -7066
rect 136422 -7622 171866 -7066
rect 172422 -7622 207866 -7066
rect 208422 -7622 243866 -7066
rect 244422 -7622 279866 -7066
rect 280422 -7622 315866 -7066
rect 316422 -7622 351866 -7066
rect 352422 -7622 387866 -7066
rect 388422 -7622 423866 -7066
rect 424422 -7622 459866 -7066
rect 460422 -7622 495866 -7066
rect 496422 -7622 531866 -7066
rect 532422 -7622 567866 -7066
rect 568422 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 0
transform 1 0 12000 0 1 3000
box 0 0 560000 349840
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 1200 0 0 0 analog_io[0]
port 1 nsew
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 560 90 0 0 analog_io[10]
port 2 nsew
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 560 90 0 0 analog_io[11]
port 3 nsew
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 560 90 0 0 analog_io[12]
port 4 nsew
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 560 90 0 0 analog_io[13]
port 5 nsew
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 560 90 0 0 analog_io[14]
port 6 nsew
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 560 90 0 0 analog_io[15]
port 7 nsew
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 560 90 0 0 analog_io[16]
port 8 nsew
flabel metal3 s -960 697220 480 697460 0 FreeSans 1200 0 0 0 analog_io[17]
port 9 nsew
flabel metal3 s -960 644996 480 645236 0 FreeSans 1200 0 0 0 analog_io[18]
port 10 nsew
flabel metal3 s -960 592908 480 593148 0 FreeSans 1200 0 0 0 analog_io[19]
port 11 nsew
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 1200 0 0 0 analog_io[1]
port 12 nsew
flabel metal3 s -960 540684 480 540924 0 FreeSans 1200 0 0 0 analog_io[20]
port 13 nsew
flabel metal3 s -960 488596 480 488836 0 FreeSans 1200 0 0 0 analog_io[21]
port 14 nsew
flabel metal3 s -960 436508 480 436748 0 FreeSans 1200 0 0 0 analog_io[22]
port 15 nsew
flabel metal3 s -960 384284 480 384524 0 FreeSans 1200 0 0 0 analog_io[23]
port 16 nsew
flabel metal3 s -960 332196 480 332436 0 FreeSans 1200 0 0 0 analog_io[24]
port 17 nsew
flabel metal3 s -960 279972 480 280212 0 FreeSans 1200 0 0 0 analog_io[25]
port 18 nsew
flabel metal3 s -960 227884 480 228124 0 FreeSans 1200 0 0 0 analog_io[26]
port 19 nsew
flabel metal3 s -960 175796 480 176036 0 FreeSans 1200 0 0 0 analog_io[27]
port 20 nsew
flabel metal3 s -960 123572 480 123812 0 FreeSans 1200 0 0 0 analog_io[28]
port 21 nsew
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 1200 0 0 0 analog_io[2]
port 22 nsew
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 1200 0 0 0 analog_io[3]
port 23 nsew
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 1200 0 0 0 analog_io[4]
port 24 nsew
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 1200 0 0 0 analog_io[5]
port 25 nsew
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 1200 0 0 0 analog_io[6]
port 26 nsew
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 1200 0 0 0 analog_io[7]
port 27 nsew
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 560 90 0 0 analog_io[8]
port 28 nsew
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 560 90 0 0 analog_io[9]
port 29 nsew
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 1200 0 0 0 io_in[0]
port 30 nsew
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 1200 0 0 0 io_in[10]
port 31 nsew
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 1200 0 0 0 io_in[11]
port 32 nsew
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 1200 0 0 0 io_in[12]
port 33 nsew
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 1200 0 0 0 io_in[13]
port 34 nsew
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 1200 0 0 0 io_in[14]
port 35 nsew
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 560 90 0 0 io_in[15]
port 36 nsew
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 560 90 0 0 io_in[16]
port 37 nsew
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 560 90 0 0 io_in[17]
port 38 nsew
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 560 90 0 0 io_in[18]
port 39 nsew
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 560 90 0 0 io_in[19]
port 40 nsew
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 1200 0 0 0 io_in[1]
port 41 nsew
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 560 90 0 0 io_in[20]
port 42 nsew
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 560 90 0 0 io_in[21]
port 43 nsew
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 560 90 0 0 io_in[22]
port 44 nsew
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 560 90 0 0 io_in[23]
port 45 nsew
flabel metal3 s -960 684164 480 684404 0 FreeSans 1200 0 0 0 io_in[24]
port 46 nsew
flabel metal3 s -960 631940 480 632180 0 FreeSans 1200 0 0 0 io_in[25]
port 47 nsew
flabel metal3 s -960 579852 480 580092 0 FreeSans 1200 0 0 0 io_in[26]
port 48 nsew
flabel metal3 s -960 527764 480 528004 0 FreeSans 1200 0 0 0 io_in[27]
port 49 nsew
flabel metal3 s -960 475540 480 475780 0 FreeSans 1200 0 0 0 io_in[28]
port 50 nsew
flabel metal3 s -960 423452 480 423692 0 FreeSans 1200 0 0 0 io_in[29]
port 51 nsew
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 1200 0 0 0 io_in[2]
port 52 nsew
flabel metal3 s -960 371228 480 371468 0 FreeSans 1200 0 0 0 io_in[30]
port 53 nsew
flabel metal3 s -960 319140 480 319380 0 FreeSans 1200 0 0 0 io_in[31]
port 54 nsew
flabel metal3 s -960 267052 480 267292 0 FreeSans 1200 0 0 0 io_in[32]
port 55 nsew
flabel metal3 s -960 214828 480 215068 0 FreeSans 1200 0 0 0 io_in[33]
port 56 nsew
flabel metal3 s -960 162740 480 162980 0 FreeSans 1200 0 0 0 io_in[34]
port 57 nsew
flabel metal3 s -960 110516 480 110756 0 FreeSans 1200 0 0 0 io_in[35]
port 58 nsew
flabel metal3 s -960 71484 480 71724 0 FreeSans 1200 0 0 0 io_in[36]
port 59 nsew
flabel metal3 s -960 32316 480 32556 0 FreeSans 1200 0 0 0 io_in[37]
port 60 nsew
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 1200 0 0 0 io_in[3]
port 61 nsew
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 1200 0 0 0 io_in[4]
port 62 nsew
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 1200 0 0 0 io_in[5]
port 63 nsew
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 1200 0 0 0 io_in[6]
port 64 nsew
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 1200 0 0 0 io_in[7]
port 65 nsew
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 1200 0 0 0 io_in[8]
port 66 nsew
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 1200 0 0 0 io_in[9]
port 67 nsew
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 1200 0 0 0 io_oeb[0]
port 68 nsew
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 1200 0 0 0 io_oeb[10]
port 69 nsew
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 1200 0 0 0 io_oeb[11]
port 70 nsew
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 1200 0 0 0 io_oeb[12]
port 71 nsew
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 1200 0 0 0 io_oeb[13]
port 72 nsew
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 1200 0 0 0 io_oeb[14]
port 73 nsew
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 560 90 0 0 io_oeb[15]
port 74 nsew
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 560 90 0 0 io_oeb[16]
port 75 nsew
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 560 90 0 0 io_oeb[17]
port 76 nsew
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 560 90 0 0 io_oeb[18]
port 77 nsew
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 560 90 0 0 io_oeb[19]
port 78 nsew
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 1200 0 0 0 io_oeb[1]
port 79 nsew
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 560 90 0 0 io_oeb[20]
port 80 nsew
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 560 90 0 0 io_oeb[21]
port 81 nsew
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 560 90 0 0 io_oeb[22]
port 82 nsew
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 560 90 0 0 io_oeb[23]
port 83 nsew
flabel metal3 s -960 658052 480 658292 0 FreeSans 1200 0 0 0 io_oeb[24]
port 84 nsew
flabel metal3 s -960 605964 480 606204 0 FreeSans 1200 0 0 0 io_oeb[25]
port 85 nsew
flabel metal3 s -960 553740 480 553980 0 FreeSans 1200 0 0 0 io_oeb[26]
port 86 nsew
flabel metal3 s -960 501652 480 501892 0 FreeSans 1200 0 0 0 io_oeb[27]
port 87 nsew
flabel metal3 s -960 449428 480 449668 0 FreeSans 1200 0 0 0 io_oeb[28]
port 88 nsew
flabel metal3 s -960 397340 480 397580 0 FreeSans 1200 0 0 0 io_oeb[29]
port 89 nsew
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 1200 0 0 0 io_oeb[2]
port 90 nsew
flabel metal3 s -960 345252 480 345492 0 FreeSans 1200 0 0 0 io_oeb[30]
port 91 nsew
flabel metal3 s -960 293028 480 293268 0 FreeSans 1200 0 0 0 io_oeb[31]
port 92 nsew
flabel metal3 s -960 240940 480 241180 0 FreeSans 1200 0 0 0 io_oeb[32]
port 93 nsew
flabel metal3 s -960 188716 480 188956 0 FreeSans 1200 0 0 0 io_oeb[33]
port 94 nsew
flabel metal3 s -960 136628 480 136868 0 FreeSans 1200 0 0 0 io_oeb[34]
port 95 nsew
flabel metal3 s -960 84540 480 84780 0 FreeSans 1200 0 0 0 io_oeb[35]
port 96 nsew
flabel metal3 s -960 45372 480 45612 0 FreeSans 1200 0 0 0 io_oeb[36]
port 97 nsew
flabel metal3 s -960 6340 480 6580 0 FreeSans 1200 0 0 0 io_oeb[37]
port 98 nsew
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 1200 0 0 0 io_oeb[3]
port 99 nsew
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 1200 0 0 0 io_oeb[4]
port 100 nsew
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 1200 0 0 0 io_oeb[5]
port 101 nsew
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 1200 0 0 0 io_oeb[6]
port 102 nsew
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 1200 0 0 0 io_oeb[7]
port 103 nsew
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 1200 0 0 0 io_oeb[8]
port 104 nsew
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 1200 0 0 0 io_oeb[9]
port 105 nsew
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 1200 0 0 0 io_out[0]
port 106 nsew
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 1200 0 0 0 io_out[10]
port 107 nsew
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 1200 0 0 0 io_out[11]
port 108 nsew
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 1200 0 0 0 io_out[12]
port 109 nsew
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 1200 0 0 0 io_out[13]
port 110 nsew
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 1200 0 0 0 io_out[14]
port 111 nsew
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 560 90 0 0 io_out[15]
port 112 nsew
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 560 90 0 0 io_out[16]
port 113 nsew
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 560 90 0 0 io_out[17]
port 114 nsew
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 560 90 0 0 io_out[18]
port 115 nsew
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 560 90 0 0 io_out[19]
port 116 nsew
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 1200 0 0 0 io_out[1]
port 117 nsew
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 560 90 0 0 io_out[20]
port 118 nsew
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 560 90 0 0 io_out[21]
port 119 nsew
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 560 90 0 0 io_out[22]
port 120 nsew
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 560 90 0 0 io_out[23]
port 121 nsew
flabel metal3 s -960 671108 480 671348 0 FreeSans 1200 0 0 0 io_out[24]
port 122 nsew
flabel metal3 s -960 619020 480 619260 0 FreeSans 1200 0 0 0 io_out[25]
port 123 nsew
flabel metal3 s -960 566796 480 567036 0 FreeSans 1200 0 0 0 io_out[26]
port 124 nsew
flabel metal3 s -960 514708 480 514948 0 FreeSans 1200 0 0 0 io_out[27]
port 125 nsew
flabel metal3 s -960 462484 480 462724 0 FreeSans 1200 0 0 0 io_out[28]
port 126 nsew
flabel metal3 s -960 410396 480 410636 0 FreeSans 1200 0 0 0 io_out[29]
port 127 nsew
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 1200 0 0 0 io_out[2]
port 128 nsew
flabel metal3 s -960 358308 480 358548 0 FreeSans 1200 0 0 0 io_out[30]
port 129 nsew
flabel metal3 s -960 306084 480 306324 0 FreeSans 1200 0 0 0 io_out[31]
port 130 nsew
flabel metal3 s -960 253996 480 254236 0 FreeSans 1200 0 0 0 io_out[32]
port 131 nsew
flabel metal3 s -960 201772 480 202012 0 FreeSans 1200 0 0 0 io_out[33]
port 132 nsew
flabel metal3 s -960 149684 480 149924 0 FreeSans 1200 0 0 0 io_out[34]
port 133 nsew
flabel metal3 s -960 97460 480 97700 0 FreeSans 1200 0 0 0 io_out[35]
port 134 nsew
flabel metal3 s -960 58428 480 58668 0 FreeSans 1200 0 0 0 io_out[36]
port 135 nsew
flabel metal3 s -960 19260 480 19500 0 FreeSans 1200 0 0 0 io_out[37]
port 136 nsew
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 1200 0 0 0 io_out[3]
port 137 nsew
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 1200 0 0 0 io_out[4]
port 138 nsew
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 1200 0 0 0 io_out[5]
port 139 nsew
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 1200 0 0 0 io_out[6]
port 140 nsew
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 1200 0 0 0 io_out[7]
port 141 nsew
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 1200 0 0 0 io_out[8]
port 142 nsew
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 1200 0 0 0 io_out[9]
port 143 nsew
flabel metal2 s 125846 -960 125958 480 0 FreeSans 560 90 0 0 la_data_in[0]
port 144 nsew
flabel metal2 s 480506 -960 480618 480 0 FreeSans 560 90 0 0 la_data_in[100]
port 145 nsew
flabel metal2 s 484002 -960 484114 480 0 FreeSans 560 90 0 0 la_data_in[101]
port 146 nsew
flabel metal2 s 487590 -960 487702 480 0 FreeSans 560 90 0 0 la_data_in[102]
port 147 nsew
flabel metal2 s 491086 -960 491198 480 0 FreeSans 560 90 0 0 la_data_in[103]
port 148 nsew
flabel metal2 s 494674 -960 494786 480 0 FreeSans 560 90 0 0 la_data_in[104]
port 149 nsew
flabel metal2 s 498170 -960 498282 480 0 FreeSans 560 90 0 0 la_data_in[105]
port 150 nsew
flabel metal2 s 501758 -960 501870 480 0 FreeSans 560 90 0 0 la_data_in[106]
port 151 nsew
flabel metal2 s 505346 -960 505458 480 0 FreeSans 560 90 0 0 la_data_in[107]
port 152 nsew
flabel metal2 s 508842 -960 508954 480 0 FreeSans 560 90 0 0 la_data_in[108]
port 153 nsew
flabel metal2 s 512430 -960 512542 480 0 FreeSans 560 90 0 0 la_data_in[109]
port 154 nsew
flabel metal2 s 161266 -960 161378 480 0 FreeSans 560 90 0 0 la_data_in[10]
port 155 nsew
flabel metal2 s 515926 -960 516038 480 0 FreeSans 560 90 0 0 la_data_in[110]
port 156 nsew
flabel metal2 s 519514 -960 519626 480 0 FreeSans 560 90 0 0 la_data_in[111]
port 157 nsew
flabel metal2 s 523010 -960 523122 480 0 FreeSans 560 90 0 0 la_data_in[112]
port 158 nsew
flabel metal2 s 526598 -960 526710 480 0 FreeSans 560 90 0 0 la_data_in[113]
port 159 nsew
flabel metal2 s 530094 -960 530206 480 0 FreeSans 560 90 0 0 la_data_in[114]
port 160 nsew
flabel metal2 s 533682 -960 533794 480 0 FreeSans 560 90 0 0 la_data_in[115]
port 161 nsew
flabel metal2 s 537178 -960 537290 480 0 FreeSans 560 90 0 0 la_data_in[116]
port 162 nsew
flabel metal2 s 540766 -960 540878 480 0 FreeSans 560 90 0 0 la_data_in[117]
port 163 nsew
flabel metal2 s 544354 -960 544466 480 0 FreeSans 560 90 0 0 la_data_in[118]
port 164 nsew
flabel metal2 s 547850 -960 547962 480 0 FreeSans 560 90 0 0 la_data_in[119]
port 165 nsew
flabel metal2 s 164854 -960 164966 480 0 FreeSans 560 90 0 0 la_data_in[11]
port 166 nsew
flabel metal2 s 551438 -960 551550 480 0 FreeSans 560 90 0 0 la_data_in[120]
port 167 nsew
flabel metal2 s 554934 -960 555046 480 0 FreeSans 560 90 0 0 la_data_in[121]
port 168 nsew
flabel metal2 s 558522 -960 558634 480 0 FreeSans 560 90 0 0 la_data_in[122]
port 169 nsew
flabel metal2 s 562018 -960 562130 480 0 FreeSans 560 90 0 0 la_data_in[123]
port 170 nsew
flabel metal2 s 565606 -960 565718 480 0 FreeSans 560 90 0 0 la_data_in[124]
port 171 nsew
flabel metal2 s 569102 -960 569214 480 0 FreeSans 560 90 0 0 la_data_in[125]
port 172 nsew
flabel metal2 s 572690 -960 572802 480 0 FreeSans 560 90 0 0 la_data_in[126]
port 173 nsew
flabel metal2 s 576278 -960 576390 480 0 FreeSans 560 90 0 0 la_data_in[127]
port 174 nsew
flabel metal2 s 168350 -960 168462 480 0 FreeSans 560 90 0 0 la_data_in[12]
port 175 nsew
flabel metal2 s 171938 -960 172050 480 0 FreeSans 560 90 0 0 la_data_in[13]
port 176 nsew
flabel metal2 s 175434 -960 175546 480 0 FreeSans 560 90 0 0 la_data_in[14]
port 177 nsew
flabel metal2 s 179022 -960 179134 480 0 FreeSans 560 90 0 0 la_data_in[15]
port 178 nsew
flabel metal2 s 182518 -960 182630 480 0 FreeSans 560 90 0 0 la_data_in[16]
port 179 nsew
flabel metal2 s 186106 -960 186218 480 0 FreeSans 560 90 0 0 la_data_in[17]
port 180 nsew
flabel metal2 s 189694 -960 189806 480 0 FreeSans 560 90 0 0 la_data_in[18]
port 181 nsew
flabel metal2 s 193190 -960 193302 480 0 FreeSans 560 90 0 0 la_data_in[19]
port 182 nsew
flabel metal2 s 129342 -960 129454 480 0 FreeSans 560 90 0 0 la_data_in[1]
port 183 nsew
flabel metal2 s 196778 -960 196890 480 0 FreeSans 560 90 0 0 la_data_in[20]
port 184 nsew
flabel metal2 s 200274 -960 200386 480 0 FreeSans 560 90 0 0 la_data_in[21]
port 185 nsew
flabel metal2 s 203862 -960 203974 480 0 FreeSans 560 90 0 0 la_data_in[22]
port 186 nsew
flabel metal2 s 207358 -960 207470 480 0 FreeSans 560 90 0 0 la_data_in[23]
port 187 nsew
flabel metal2 s 210946 -960 211058 480 0 FreeSans 560 90 0 0 la_data_in[24]
port 188 nsew
flabel metal2 s 214442 -960 214554 480 0 FreeSans 560 90 0 0 la_data_in[25]
port 189 nsew
flabel metal2 s 218030 -960 218142 480 0 FreeSans 560 90 0 0 la_data_in[26]
port 190 nsew
flabel metal2 s 221526 -960 221638 480 0 FreeSans 560 90 0 0 la_data_in[27]
port 191 nsew
flabel metal2 s 225114 -960 225226 480 0 FreeSans 560 90 0 0 la_data_in[28]
port 192 nsew
flabel metal2 s 228702 -960 228814 480 0 FreeSans 560 90 0 0 la_data_in[29]
port 193 nsew
flabel metal2 s 132930 -960 133042 480 0 FreeSans 560 90 0 0 la_data_in[2]
port 194 nsew
flabel metal2 s 232198 -960 232310 480 0 FreeSans 560 90 0 0 la_data_in[30]
port 195 nsew
flabel metal2 s 235786 -960 235898 480 0 FreeSans 560 90 0 0 la_data_in[31]
port 196 nsew
flabel metal2 s 239282 -960 239394 480 0 FreeSans 560 90 0 0 la_data_in[32]
port 197 nsew
flabel metal2 s 242870 -960 242982 480 0 FreeSans 560 90 0 0 la_data_in[33]
port 198 nsew
flabel metal2 s 246366 -960 246478 480 0 FreeSans 560 90 0 0 la_data_in[34]
port 199 nsew
flabel metal2 s 249954 -960 250066 480 0 FreeSans 560 90 0 0 la_data_in[35]
port 200 nsew
flabel metal2 s 253450 -960 253562 480 0 FreeSans 560 90 0 0 la_data_in[36]
port 201 nsew
flabel metal2 s 257038 -960 257150 480 0 FreeSans 560 90 0 0 la_data_in[37]
port 202 nsew
flabel metal2 s 260626 -960 260738 480 0 FreeSans 560 90 0 0 la_data_in[38]
port 203 nsew
flabel metal2 s 264122 -960 264234 480 0 FreeSans 560 90 0 0 la_data_in[39]
port 204 nsew
flabel metal2 s 136426 -960 136538 480 0 FreeSans 560 90 0 0 la_data_in[3]
port 205 nsew
flabel metal2 s 267710 -960 267822 480 0 FreeSans 560 90 0 0 la_data_in[40]
port 206 nsew
flabel metal2 s 271206 -960 271318 480 0 FreeSans 560 90 0 0 la_data_in[41]
port 207 nsew
flabel metal2 s 274794 -960 274906 480 0 FreeSans 560 90 0 0 la_data_in[42]
port 208 nsew
flabel metal2 s 278290 -960 278402 480 0 FreeSans 560 90 0 0 la_data_in[43]
port 209 nsew
flabel metal2 s 281878 -960 281990 480 0 FreeSans 560 90 0 0 la_data_in[44]
port 210 nsew
flabel metal2 s 285374 -960 285486 480 0 FreeSans 560 90 0 0 la_data_in[45]
port 211 nsew
flabel metal2 s 288962 -960 289074 480 0 FreeSans 560 90 0 0 la_data_in[46]
port 212 nsew
flabel metal2 s 292550 -960 292662 480 0 FreeSans 560 90 0 0 la_data_in[47]
port 213 nsew
flabel metal2 s 296046 -960 296158 480 0 FreeSans 560 90 0 0 la_data_in[48]
port 214 nsew
flabel metal2 s 299634 -960 299746 480 0 FreeSans 560 90 0 0 la_data_in[49]
port 215 nsew
flabel metal2 s 140014 -960 140126 480 0 FreeSans 560 90 0 0 la_data_in[4]
port 216 nsew
flabel metal2 s 303130 -960 303242 480 0 FreeSans 560 90 0 0 la_data_in[50]
port 217 nsew
flabel metal2 s 306718 -960 306830 480 0 FreeSans 560 90 0 0 la_data_in[51]
port 218 nsew
flabel metal2 s 310214 -960 310326 480 0 FreeSans 560 90 0 0 la_data_in[52]
port 219 nsew
flabel metal2 s 313802 -960 313914 480 0 FreeSans 560 90 0 0 la_data_in[53]
port 220 nsew
flabel metal2 s 317298 -960 317410 480 0 FreeSans 560 90 0 0 la_data_in[54]
port 221 nsew
flabel metal2 s 320886 -960 320998 480 0 FreeSans 560 90 0 0 la_data_in[55]
port 222 nsew
flabel metal2 s 324382 -960 324494 480 0 FreeSans 560 90 0 0 la_data_in[56]
port 223 nsew
flabel metal2 s 327970 -960 328082 480 0 FreeSans 560 90 0 0 la_data_in[57]
port 224 nsew
flabel metal2 s 331558 -960 331670 480 0 FreeSans 560 90 0 0 la_data_in[58]
port 225 nsew
flabel metal2 s 335054 -960 335166 480 0 FreeSans 560 90 0 0 la_data_in[59]
port 226 nsew
flabel metal2 s 143510 -960 143622 480 0 FreeSans 560 90 0 0 la_data_in[5]
port 227 nsew
flabel metal2 s 338642 -960 338754 480 0 FreeSans 560 90 0 0 la_data_in[60]
port 228 nsew
flabel metal2 s 342138 -960 342250 480 0 FreeSans 560 90 0 0 la_data_in[61]
port 229 nsew
flabel metal2 s 345726 -960 345838 480 0 FreeSans 560 90 0 0 la_data_in[62]
port 230 nsew
flabel metal2 s 349222 -960 349334 480 0 FreeSans 560 90 0 0 la_data_in[63]
port 231 nsew
flabel metal2 s 352810 -960 352922 480 0 FreeSans 560 90 0 0 la_data_in[64]
port 232 nsew
flabel metal2 s 356306 -960 356418 480 0 FreeSans 560 90 0 0 la_data_in[65]
port 233 nsew
flabel metal2 s 359894 -960 360006 480 0 FreeSans 560 90 0 0 la_data_in[66]
port 234 nsew
flabel metal2 s 363482 -960 363594 480 0 FreeSans 560 90 0 0 la_data_in[67]
port 235 nsew
flabel metal2 s 366978 -960 367090 480 0 FreeSans 560 90 0 0 la_data_in[68]
port 236 nsew
flabel metal2 s 370566 -960 370678 480 0 FreeSans 560 90 0 0 la_data_in[69]
port 237 nsew
flabel metal2 s 147098 -960 147210 480 0 FreeSans 560 90 0 0 la_data_in[6]
port 238 nsew
flabel metal2 s 374062 -960 374174 480 0 FreeSans 560 90 0 0 la_data_in[70]
port 239 nsew
flabel metal2 s 377650 -960 377762 480 0 FreeSans 560 90 0 0 la_data_in[71]
port 240 nsew
flabel metal2 s 381146 -960 381258 480 0 FreeSans 560 90 0 0 la_data_in[72]
port 241 nsew
flabel metal2 s 384734 -960 384846 480 0 FreeSans 560 90 0 0 la_data_in[73]
port 242 nsew
flabel metal2 s 388230 -960 388342 480 0 FreeSans 560 90 0 0 la_data_in[74]
port 243 nsew
flabel metal2 s 391818 -960 391930 480 0 FreeSans 560 90 0 0 la_data_in[75]
port 244 nsew
flabel metal2 s 395314 -960 395426 480 0 FreeSans 560 90 0 0 la_data_in[76]
port 245 nsew
flabel metal2 s 398902 -960 399014 480 0 FreeSans 560 90 0 0 la_data_in[77]
port 246 nsew
flabel metal2 s 402490 -960 402602 480 0 FreeSans 560 90 0 0 la_data_in[78]
port 247 nsew
flabel metal2 s 405986 -960 406098 480 0 FreeSans 560 90 0 0 la_data_in[79]
port 248 nsew
flabel metal2 s 150594 -960 150706 480 0 FreeSans 560 90 0 0 la_data_in[7]
port 249 nsew
flabel metal2 s 409574 -960 409686 480 0 FreeSans 560 90 0 0 la_data_in[80]
port 250 nsew
flabel metal2 s 413070 -960 413182 480 0 FreeSans 560 90 0 0 la_data_in[81]
port 251 nsew
flabel metal2 s 416658 -960 416770 480 0 FreeSans 560 90 0 0 la_data_in[82]
port 252 nsew
flabel metal2 s 420154 -960 420266 480 0 FreeSans 560 90 0 0 la_data_in[83]
port 253 nsew
flabel metal2 s 423742 -960 423854 480 0 FreeSans 560 90 0 0 la_data_in[84]
port 254 nsew
flabel metal2 s 427238 -960 427350 480 0 FreeSans 560 90 0 0 la_data_in[85]
port 255 nsew
flabel metal2 s 430826 -960 430938 480 0 FreeSans 560 90 0 0 la_data_in[86]
port 256 nsew
flabel metal2 s 434414 -960 434526 480 0 FreeSans 560 90 0 0 la_data_in[87]
port 257 nsew
flabel metal2 s 437910 -960 438022 480 0 FreeSans 560 90 0 0 la_data_in[88]
port 258 nsew
flabel metal2 s 441498 -960 441610 480 0 FreeSans 560 90 0 0 la_data_in[89]
port 259 nsew
flabel metal2 s 154182 -960 154294 480 0 FreeSans 560 90 0 0 la_data_in[8]
port 260 nsew
flabel metal2 s 444994 -960 445106 480 0 FreeSans 560 90 0 0 la_data_in[90]
port 261 nsew
flabel metal2 s 448582 -960 448694 480 0 FreeSans 560 90 0 0 la_data_in[91]
port 262 nsew
flabel metal2 s 452078 -960 452190 480 0 FreeSans 560 90 0 0 la_data_in[92]
port 263 nsew
flabel metal2 s 455666 -960 455778 480 0 FreeSans 560 90 0 0 la_data_in[93]
port 264 nsew
flabel metal2 s 459162 -960 459274 480 0 FreeSans 560 90 0 0 la_data_in[94]
port 265 nsew
flabel metal2 s 462750 -960 462862 480 0 FreeSans 560 90 0 0 la_data_in[95]
port 266 nsew
flabel metal2 s 466246 -960 466358 480 0 FreeSans 560 90 0 0 la_data_in[96]
port 267 nsew
flabel metal2 s 469834 -960 469946 480 0 FreeSans 560 90 0 0 la_data_in[97]
port 268 nsew
flabel metal2 s 473422 -960 473534 480 0 FreeSans 560 90 0 0 la_data_in[98]
port 269 nsew
flabel metal2 s 476918 -960 477030 480 0 FreeSans 560 90 0 0 la_data_in[99]
port 270 nsew
flabel metal2 s 157770 -960 157882 480 0 FreeSans 560 90 0 0 la_data_in[9]
port 271 nsew
flabel metal2 s 126950 -960 127062 480 0 FreeSans 560 90 0 0 la_data_out[0]
port 272 nsew
flabel metal2 s 481702 -960 481814 480 0 FreeSans 560 90 0 0 la_data_out[100]
port 273 nsew
flabel metal2 s 485198 -960 485310 480 0 FreeSans 560 90 0 0 la_data_out[101]
port 274 nsew
flabel metal2 s 488786 -960 488898 480 0 FreeSans 560 90 0 0 la_data_out[102]
port 275 nsew
flabel metal2 s 492282 -960 492394 480 0 FreeSans 560 90 0 0 la_data_out[103]
port 276 nsew
flabel metal2 s 495870 -960 495982 480 0 FreeSans 560 90 0 0 la_data_out[104]
port 277 nsew
flabel metal2 s 499366 -960 499478 480 0 FreeSans 560 90 0 0 la_data_out[105]
port 278 nsew
flabel metal2 s 502954 -960 503066 480 0 FreeSans 560 90 0 0 la_data_out[106]
port 279 nsew
flabel metal2 s 506450 -960 506562 480 0 FreeSans 560 90 0 0 la_data_out[107]
port 280 nsew
flabel metal2 s 510038 -960 510150 480 0 FreeSans 560 90 0 0 la_data_out[108]
port 281 nsew
flabel metal2 s 513534 -960 513646 480 0 FreeSans 560 90 0 0 la_data_out[109]
port 282 nsew
flabel metal2 s 162462 -960 162574 480 0 FreeSans 560 90 0 0 la_data_out[10]
port 283 nsew
flabel metal2 s 517122 -960 517234 480 0 FreeSans 560 90 0 0 la_data_out[110]
port 284 nsew
flabel metal2 s 520710 -960 520822 480 0 FreeSans 560 90 0 0 la_data_out[111]
port 285 nsew
flabel metal2 s 524206 -960 524318 480 0 FreeSans 560 90 0 0 la_data_out[112]
port 286 nsew
flabel metal2 s 527794 -960 527906 480 0 FreeSans 560 90 0 0 la_data_out[113]
port 287 nsew
flabel metal2 s 531290 -960 531402 480 0 FreeSans 560 90 0 0 la_data_out[114]
port 288 nsew
flabel metal2 s 534878 -960 534990 480 0 FreeSans 560 90 0 0 la_data_out[115]
port 289 nsew
flabel metal2 s 538374 -960 538486 480 0 FreeSans 560 90 0 0 la_data_out[116]
port 290 nsew
flabel metal2 s 541962 -960 542074 480 0 FreeSans 560 90 0 0 la_data_out[117]
port 291 nsew
flabel metal2 s 545458 -960 545570 480 0 FreeSans 560 90 0 0 la_data_out[118]
port 292 nsew
flabel metal2 s 549046 -960 549158 480 0 FreeSans 560 90 0 0 la_data_out[119]
port 293 nsew
flabel metal2 s 166050 -960 166162 480 0 FreeSans 560 90 0 0 la_data_out[11]
port 294 nsew
flabel metal2 s 552634 -960 552746 480 0 FreeSans 560 90 0 0 la_data_out[120]
port 295 nsew
flabel metal2 s 556130 -960 556242 480 0 FreeSans 560 90 0 0 la_data_out[121]
port 296 nsew
flabel metal2 s 559718 -960 559830 480 0 FreeSans 560 90 0 0 la_data_out[122]
port 297 nsew
flabel metal2 s 563214 -960 563326 480 0 FreeSans 560 90 0 0 la_data_out[123]
port 298 nsew
flabel metal2 s 566802 -960 566914 480 0 FreeSans 560 90 0 0 la_data_out[124]
port 299 nsew
flabel metal2 s 570298 -960 570410 480 0 FreeSans 560 90 0 0 la_data_out[125]
port 300 nsew
flabel metal2 s 573886 -960 573998 480 0 FreeSans 560 90 0 0 la_data_out[126]
port 301 nsew
flabel metal2 s 577382 -960 577494 480 0 FreeSans 560 90 0 0 la_data_out[127]
port 302 nsew
flabel metal2 s 169546 -960 169658 480 0 FreeSans 560 90 0 0 la_data_out[12]
port 303 nsew
flabel metal2 s 173134 -960 173246 480 0 FreeSans 560 90 0 0 la_data_out[13]
port 304 nsew
flabel metal2 s 176630 -960 176742 480 0 FreeSans 560 90 0 0 la_data_out[14]
port 305 nsew
flabel metal2 s 180218 -960 180330 480 0 FreeSans 560 90 0 0 la_data_out[15]
port 306 nsew
flabel metal2 s 183714 -960 183826 480 0 FreeSans 560 90 0 0 la_data_out[16]
port 307 nsew
flabel metal2 s 187302 -960 187414 480 0 FreeSans 560 90 0 0 la_data_out[17]
port 308 nsew
flabel metal2 s 190798 -960 190910 480 0 FreeSans 560 90 0 0 la_data_out[18]
port 309 nsew
flabel metal2 s 194386 -960 194498 480 0 FreeSans 560 90 0 0 la_data_out[19]
port 310 nsew
flabel metal2 s 130538 -960 130650 480 0 FreeSans 560 90 0 0 la_data_out[1]
port 311 nsew
flabel metal2 s 197882 -960 197994 480 0 FreeSans 560 90 0 0 la_data_out[20]
port 312 nsew
flabel metal2 s 201470 -960 201582 480 0 FreeSans 560 90 0 0 la_data_out[21]
port 313 nsew
flabel metal2 s 205058 -960 205170 480 0 FreeSans 560 90 0 0 la_data_out[22]
port 314 nsew
flabel metal2 s 208554 -960 208666 480 0 FreeSans 560 90 0 0 la_data_out[23]
port 315 nsew
flabel metal2 s 212142 -960 212254 480 0 FreeSans 560 90 0 0 la_data_out[24]
port 316 nsew
flabel metal2 s 215638 -960 215750 480 0 FreeSans 560 90 0 0 la_data_out[25]
port 317 nsew
flabel metal2 s 219226 -960 219338 480 0 FreeSans 560 90 0 0 la_data_out[26]
port 318 nsew
flabel metal2 s 222722 -960 222834 480 0 FreeSans 560 90 0 0 la_data_out[27]
port 319 nsew
flabel metal2 s 226310 -960 226422 480 0 FreeSans 560 90 0 0 la_data_out[28]
port 320 nsew
flabel metal2 s 229806 -960 229918 480 0 FreeSans 560 90 0 0 la_data_out[29]
port 321 nsew
flabel metal2 s 134126 -960 134238 480 0 FreeSans 560 90 0 0 la_data_out[2]
port 322 nsew
flabel metal2 s 233394 -960 233506 480 0 FreeSans 560 90 0 0 la_data_out[30]
port 323 nsew
flabel metal2 s 236982 -960 237094 480 0 FreeSans 560 90 0 0 la_data_out[31]
port 324 nsew
flabel metal2 s 240478 -960 240590 480 0 FreeSans 560 90 0 0 la_data_out[32]
port 325 nsew
flabel metal2 s 244066 -960 244178 480 0 FreeSans 560 90 0 0 la_data_out[33]
port 326 nsew
flabel metal2 s 247562 -960 247674 480 0 FreeSans 560 90 0 0 la_data_out[34]
port 327 nsew
flabel metal2 s 251150 -960 251262 480 0 FreeSans 560 90 0 0 la_data_out[35]
port 328 nsew
flabel metal2 s 254646 -960 254758 480 0 FreeSans 560 90 0 0 la_data_out[36]
port 329 nsew
flabel metal2 s 258234 -960 258346 480 0 FreeSans 560 90 0 0 la_data_out[37]
port 330 nsew
flabel metal2 s 261730 -960 261842 480 0 FreeSans 560 90 0 0 la_data_out[38]
port 331 nsew
flabel metal2 s 265318 -960 265430 480 0 FreeSans 560 90 0 0 la_data_out[39]
port 332 nsew
flabel metal2 s 137622 -960 137734 480 0 FreeSans 560 90 0 0 la_data_out[3]
port 333 nsew
flabel metal2 s 268814 -960 268926 480 0 FreeSans 560 90 0 0 la_data_out[40]
port 334 nsew
flabel metal2 s 272402 -960 272514 480 0 FreeSans 560 90 0 0 la_data_out[41]
port 335 nsew
flabel metal2 s 275990 -960 276102 480 0 FreeSans 560 90 0 0 la_data_out[42]
port 336 nsew
flabel metal2 s 279486 -960 279598 480 0 FreeSans 560 90 0 0 la_data_out[43]
port 337 nsew
flabel metal2 s 283074 -960 283186 480 0 FreeSans 560 90 0 0 la_data_out[44]
port 338 nsew
flabel metal2 s 286570 -960 286682 480 0 FreeSans 560 90 0 0 la_data_out[45]
port 339 nsew
flabel metal2 s 290158 -960 290270 480 0 FreeSans 560 90 0 0 la_data_out[46]
port 340 nsew
flabel metal2 s 293654 -960 293766 480 0 FreeSans 560 90 0 0 la_data_out[47]
port 341 nsew
flabel metal2 s 297242 -960 297354 480 0 FreeSans 560 90 0 0 la_data_out[48]
port 342 nsew
flabel metal2 s 300738 -960 300850 480 0 FreeSans 560 90 0 0 la_data_out[49]
port 343 nsew
flabel metal2 s 141210 -960 141322 480 0 FreeSans 560 90 0 0 la_data_out[4]
port 344 nsew
flabel metal2 s 304326 -960 304438 480 0 FreeSans 560 90 0 0 la_data_out[50]
port 345 nsew
flabel metal2 s 307914 -960 308026 480 0 FreeSans 560 90 0 0 la_data_out[51]
port 346 nsew
flabel metal2 s 311410 -960 311522 480 0 FreeSans 560 90 0 0 la_data_out[52]
port 347 nsew
flabel metal2 s 314998 -960 315110 480 0 FreeSans 560 90 0 0 la_data_out[53]
port 348 nsew
flabel metal2 s 318494 -960 318606 480 0 FreeSans 560 90 0 0 la_data_out[54]
port 349 nsew
flabel metal2 s 322082 -960 322194 480 0 FreeSans 560 90 0 0 la_data_out[55]
port 350 nsew
flabel metal2 s 325578 -960 325690 480 0 FreeSans 560 90 0 0 la_data_out[56]
port 351 nsew
flabel metal2 s 329166 -960 329278 480 0 FreeSans 560 90 0 0 la_data_out[57]
port 352 nsew
flabel metal2 s 332662 -960 332774 480 0 FreeSans 560 90 0 0 la_data_out[58]
port 353 nsew
flabel metal2 s 336250 -960 336362 480 0 FreeSans 560 90 0 0 la_data_out[59]
port 354 nsew
flabel metal2 s 144706 -960 144818 480 0 FreeSans 560 90 0 0 la_data_out[5]
port 355 nsew
flabel metal2 s 339838 -960 339950 480 0 FreeSans 560 90 0 0 la_data_out[60]
port 356 nsew
flabel metal2 s 343334 -960 343446 480 0 FreeSans 560 90 0 0 la_data_out[61]
port 357 nsew
flabel metal2 s 346922 -960 347034 480 0 FreeSans 560 90 0 0 la_data_out[62]
port 358 nsew
flabel metal2 s 350418 -960 350530 480 0 FreeSans 560 90 0 0 la_data_out[63]
port 359 nsew
flabel metal2 s 354006 -960 354118 480 0 FreeSans 560 90 0 0 la_data_out[64]
port 360 nsew
flabel metal2 s 357502 -960 357614 480 0 FreeSans 560 90 0 0 la_data_out[65]
port 361 nsew
flabel metal2 s 361090 -960 361202 480 0 FreeSans 560 90 0 0 la_data_out[66]
port 362 nsew
flabel metal2 s 364586 -960 364698 480 0 FreeSans 560 90 0 0 la_data_out[67]
port 363 nsew
flabel metal2 s 368174 -960 368286 480 0 FreeSans 560 90 0 0 la_data_out[68]
port 364 nsew
flabel metal2 s 371670 -960 371782 480 0 FreeSans 560 90 0 0 la_data_out[69]
port 365 nsew
flabel metal2 s 148294 -960 148406 480 0 FreeSans 560 90 0 0 la_data_out[6]
port 366 nsew
flabel metal2 s 375258 -960 375370 480 0 FreeSans 560 90 0 0 la_data_out[70]
port 367 nsew
flabel metal2 s 378846 -960 378958 480 0 FreeSans 560 90 0 0 la_data_out[71]
port 368 nsew
flabel metal2 s 382342 -960 382454 480 0 FreeSans 560 90 0 0 la_data_out[72]
port 369 nsew
flabel metal2 s 385930 -960 386042 480 0 FreeSans 560 90 0 0 la_data_out[73]
port 370 nsew
flabel metal2 s 389426 -960 389538 480 0 FreeSans 560 90 0 0 la_data_out[74]
port 371 nsew
flabel metal2 s 393014 -960 393126 480 0 FreeSans 560 90 0 0 la_data_out[75]
port 372 nsew
flabel metal2 s 396510 -960 396622 480 0 FreeSans 560 90 0 0 la_data_out[76]
port 373 nsew
flabel metal2 s 400098 -960 400210 480 0 FreeSans 560 90 0 0 la_data_out[77]
port 374 nsew
flabel metal2 s 403594 -960 403706 480 0 FreeSans 560 90 0 0 la_data_out[78]
port 375 nsew
flabel metal2 s 407182 -960 407294 480 0 FreeSans 560 90 0 0 la_data_out[79]
port 376 nsew
flabel metal2 s 151790 -960 151902 480 0 FreeSans 560 90 0 0 la_data_out[7]
port 377 nsew
flabel metal2 s 410770 -960 410882 480 0 FreeSans 560 90 0 0 la_data_out[80]
port 378 nsew
flabel metal2 s 414266 -960 414378 480 0 FreeSans 560 90 0 0 la_data_out[81]
port 379 nsew
flabel metal2 s 417854 -960 417966 480 0 FreeSans 560 90 0 0 la_data_out[82]
port 380 nsew
flabel metal2 s 421350 -960 421462 480 0 FreeSans 560 90 0 0 la_data_out[83]
port 381 nsew
flabel metal2 s 424938 -960 425050 480 0 FreeSans 560 90 0 0 la_data_out[84]
port 382 nsew
flabel metal2 s 428434 -960 428546 480 0 FreeSans 560 90 0 0 la_data_out[85]
port 383 nsew
flabel metal2 s 432022 -960 432134 480 0 FreeSans 560 90 0 0 la_data_out[86]
port 384 nsew
flabel metal2 s 435518 -960 435630 480 0 FreeSans 560 90 0 0 la_data_out[87]
port 385 nsew
flabel metal2 s 439106 -960 439218 480 0 FreeSans 560 90 0 0 la_data_out[88]
port 386 nsew
flabel metal2 s 442602 -960 442714 480 0 FreeSans 560 90 0 0 la_data_out[89]
port 387 nsew
flabel metal2 s 155378 -960 155490 480 0 FreeSans 560 90 0 0 la_data_out[8]
port 388 nsew
flabel metal2 s 446190 -960 446302 480 0 FreeSans 560 90 0 0 la_data_out[90]
port 389 nsew
flabel metal2 s 449778 -960 449890 480 0 FreeSans 560 90 0 0 la_data_out[91]
port 390 nsew
flabel metal2 s 453274 -960 453386 480 0 FreeSans 560 90 0 0 la_data_out[92]
port 391 nsew
flabel metal2 s 456862 -960 456974 480 0 FreeSans 560 90 0 0 la_data_out[93]
port 392 nsew
flabel metal2 s 460358 -960 460470 480 0 FreeSans 560 90 0 0 la_data_out[94]
port 393 nsew
flabel metal2 s 463946 -960 464058 480 0 FreeSans 560 90 0 0 la_data_out[95]
port 394 nsew
flabel metal2 s 467442 -960 467554 480 0 FreeSans 560 90 0 0 la_data_out[96]
port 395 nsew
flabel metal2 s 471030 -960 471142 480 0 FreeSans 560 90 0 0 la_data_out[97]
port 396 nsew
flabel metal2 s 474526 -960 474638 480 0 FreeSans 560 90 0 0 la_data_out[98]
port 397 nsew
flabel metal2 s 478114 -960 478226 480 0 FreeSans 560 90 0 0 la_data_out[99]
port 398 nsew
flabel metal2 s 158874 -960 158986 480 0 FreeSans 560 90 0 0 la_data_out[9]
port 399 nsew
flabel metal2 s 128146 -960 128258 480 0 FreeSans 560 90 0 0 la_oenb[0]
port 400 nsew
flabel metal2 s 482806 -960 482918 480 0 FreeSans 560 90 0 0 la_oenb[100]
port 401 nsew
flabel metal2 s 486394 -960 486506 480 0 FreeSans 560 90 0 0 la_oenb[101]
port 402 nsew
flabel metal2 s 489890 -960 490002 480 0 FreeSans 560 90 0 0 la_oenb[102]
port 403 nsew
flabel metal2 s 493478 -960 493590 480 0 FreeSans 560 90 0 0 la_oenb[103]
port 404 nsew
flabel metal2 s 497066 -960 497178 480 0 FreeSans 560 90 0 0 la_oenb[104]
port 405 nsew
flabel metal2 s 500562 -960 500674 480 0 FreeSans 560 90 0 0 la_oenb[105]
port 406 nsew
flabel metal2 s 504150 -960 504262 480 0 FreeSans 560 90 0 0 la_oenb[106]
port 407 nsew
flabel metal2 s 507646 -960 507758 480 0 FreeSans 560 90 0 0 la_oenb[107]
port 408 nsew
flabel metal2 s 511234 -960 511346 480 0 FreeSans 560 90 0 0 la_oenb[108]
port 409 nsew
flabel metal2 s 514730 -960 514842 480 0 FreeSans 560 90 0 0 la_oenb[109]
port 410 nsew
flabel metal2 s 163658 -960 163770 480 0 FreeSans 560 90 0 0 la_oenb[10]
port 411 nsew
flabel metal2 s 518318 -960 518430 480 0 FreeSans 560 90 0 0 la_oenb[110]
port 412 nsew
flabel metal2 s 521814 -960 521926 480 0 FreeSans 560 90 0 0 la_oenb[111]
port 413 nsew
flabel metal2 s 525402 -960 525514 480 0 FreeSans 560 90 0 0 la_oenb[112]
port 414 nsew
flabel metal2 s 528990 -960 529102 480 0 FreeSans 560 90 0 0 la_oenb[113]
port 415 nsew
flabel metal2 s 532486 -960 532598 480 0 FreeSans 560 90 0 0 la_oenb[114]
port 416 nsew
flabel metal2 s 536074 -960 536186 480 0 FreeSans 560 90 0 0 la_oenb[115]
port 417 nsew
flabel metal2 s 539570 -960 539682 480 0 FreeSans 560 90 0 0 la_oenb[116]
port 418 nsew
flabel metal2 s 543158 -960 543270 480 0 FreeSans 560 90 0 0 la_oenb[117]
port 419 nsew
flabel metal2 s 546654 -960 546766 480 0 FreeSans 560 90 0 0 la_oenb[118]
port 420 nsew
flabel metal2 s 550242 -960 550354 480 0 FreeSans 560 90 0 0 la_oenb[119]
port 421 nsew
flabel metal2 s 167154 -960 167266 480 0 FreeSans 560 90 0 0 la_oenb[11]
port 422 nsew
flabel metal2 s 553738 -960 553850 480 0 FreeSans 560 90 0 0 la_oenb[120]
port 423 nsew
flabel metal2 s 557326 -960 557438 480 0 FreeSans 560 90 0 0 la_oenb[121]
port 424 nsew
flabel metal2 s 560822 -960 560934 480 0 FreeSans 560 90 0 0 la_oenb[122]
port 425 nsew
flabel metal2 s 564410 -960 564522 480 0 FreeSans 560 90 0 0 la_oenb[123]
port 426 nsew
flabel metal2 s 567998 -960 568110 480 0 FreeSans 560 90 0 0 la_oenb[124]
port 427 nsew
flabel metal2 s 571494 -960 571606 480 0 FreeSans 560 90 0 0 la_oenb[125]
port 428 nsew
flabel metal2 s 575082 -960 575194 480 0 FreeSans 560 90 0 0 la_oenb[126]
port 429 nsew
flabel metal2 s 578578 -960 578690 480 0 FreeSans 560 90 0 0 la_oenb[127]
port 430 nsew
flabel metal2 s 170742 -960 170854 480 0 FreeSans 560 90 0 0 la_oenb[12]
port 431 nsew
flabel metal2 s 174238 -960 174350 480 0 FreeSans 560 90 0 0 la_oenb[13]
port 432 nsew
flabel metal2 s 177826 -960 177938 480 0 FreeSans 560 90 0 0 la_oenb[14]
port 433 nsew
flabel metal2 s 181414 -960 181526 480 0 FreeSans 560 90 0 0 la_oenb[15]
port 434 nsew
flabel metal2 s 184910 -960 185022 480 0 FreeSans 560 90 0 0 la_oenb[16]
port 435 nsew
flabel metal2 s 188498 -960 188610 480 0 FreeSans 560 90 0 0 la_oenb[17]
port 436 nsew
flabel metal2 s 191994 -960 192106 480 0 FreeSans 560 90 0 0 la_oenb[18]
port 437 nsew
flabel metal2 s 195582 -960 195694 480 0 FreeSans 560 90 0 0 la_oenb[19]
port 438 nsew
flabel metal2 s 131734 -960 131846 480 0 FreeSans 560 90 0 0 la_oenb[1]
port 439 nsew
flabel metal2 s 199078 -960 199190 480 0 FreeSans 560 90 0 0 la_oenb[20]
port 440 nsew
flabel metal2 s 202666 -960 202778 480 0 FreeSans 560 90 0 0 la_oenb[21]
port 441 nsew
flabel metal2 s 206162 -960 206274 480 0 FreeSans 560 90 0 0 la_oenb[22]
port 442 nsew
flabel metal2 s 209750 -960 209862 480 0 FreeSans 560 90 0 0 la_oenb[23]
port 443 nsew
flabel metal2 s 213338 -960 213450 480 0 FreeSans 560 90 0 0 la_oenb[24]
port 444 nsew
flabel metal2 s 216834 -960 216946 480 0 FreeSans 560 90 0 0 la_oenb[25]
port 445 nsew
flabel metal2 s 220422 -960 220534 480 0 FreeSans 560 90 0 0 la_oenb[26]
port 446 nsew
flabel metal2 s 223918 -960 224030 480 0 FreeSans 560 90 0 0 la_oenb[27]
port 447 nsew
flabel metal2 s 227506 -960 227618 480 0 FreeSans 560 90 0 0 la_oenb[28]
port 448 nsew
flabel metal2 s 231002 -960 231114 480 0 FreeSans 560 90 0 0 la_oenb[29]
port 449 nsew
flabel metal2 s 135230 -960 135342 480 0 FreeSans 560 90 0 0 la_oenb[2]
port 450 nsew
flabel metal2 s 234590 -960 234702 480 0 FreeSans 560 90 0 0 la_oenb[30]
port 451 nsew
flabel metal2 s 238086 -960 238198 480 0 FreeSans 560 90 0 0 la_oenb[31]
port 452 nsew
flabel metal2 s 241674 -960 241786 480 0 FreeSans 560 90 0 0 la_oenb[32]
port 453 nsew
flabel metal2 s 245170 -960 245282 480 0 FreeSans 560 90 0 0 la_oenb[33]
port 454 nsew
flabel metal2 s 248758 -960 248870 480 0 FreeSans 560 90 0 0 la_oenb[34]
port 455 nsew
flabel metal2 s 252346 -960 252458 480 0 FreeSans 560 90 0 0 la_oenb[35]
port 456 nsew
flabel metal2 s 255842 -960 255954 480 0 FreeSans 560 90 0 0 la_oenb[36]
port 457 nsew
flabel metal2 s 259430 -960 259542 480 0 FreeSans 560 90 0 0 la_oenb[37]
port 458 nsew
flabel metal2 s 262926 -960 263038 480 0 FreeSans 560 90 0 0 la_oenb[38]
port 459 nsew
flabel metal2 s 266514 -960 266626 480 0 FreeSans 560 90 0 0 la_oenb[39]
port 460 nsew
flabel metal2 s 138818 -960 138930 480 0 FreeSans 560 90 0 0 la_oenb[3]
port 461 nsew
flabel metal2 s 270010 -960 270122 480 0 FreeSans 560 90 0 0 la_oenb[40]
port 462 nsew
flabel metal2 s 273598 -960 273710 480 0 FreeSans 560 90 0 0 la_oenb[41]
port 463 nsew
flabel metal2 s 277094 -960 277206 480 0 FreeSans 560 90 0 0 la_oenb[42]
port 464 nsew
flabel metal2 s 280682 -960 280794 480 0 FreeSans 560 90 0 0 la_oenb[43]
port 465 nsew
flabel metal2 s 284270 -960 284382 480 0 FreeSans 560 90 0 0 la_oenb[44]
port 466 nsew
flabel metal2 s 287766 -960 287878 480 0 FreeSans 560 90 0 0 la_oenb[45]
port 467 nsew
flabel metal2 s 291354 -960 291466 480 0 FreeSans 560 90 0 0 la_oenb[46]
port 468 nsew
flabel metal2 s 294850 -960 294962 480 0 FreeSans 560 90 0 0 la_oenb[47]
port 469 nsew
flabel metal2 s 298438 -960 298550 480 0 FreeSans 560 90 0 0 la_oenb[48]
port 470 nsew
flabel metal2 s 301934 -960 302046 480 0 FreeSans 560 90 0 0 la_oenb[49]
port 471 nsew
flabel metal2 s 142406 -960 142518 480 0 FreeSans 560 90 0 0 la_oenb[4]
port 472 nsew
flabel metal2 s 305522 -960 305634 480 0 FreeSans 560 90 0 0 la_oenb[50]
port 473 nsew
flabel metal2 s 309018 -960 309130 480 0 FreeSans 560 90 0 0 la_oenb[51]
port 474 nsew
flabel metal2 s 312606 -960 312718 480 0 FreeSans 560 90 0 0 la_oenb[52]
port 475 nsew
flabel metal2 s 316194 -960 316306 480 0 FreeSans 560 90 0 0 la_oenb[53]
port 476 nsew
flabel metal2 s 319690 -960 319802 480 0 FreeSans 560 90 0 0 la_oenb[54]
port 477 nsew
flabel metal2 s 323278 -960 323390 480 0 FreeSans 560 90 0 0 la_oenb[55]
port 478 nsew
flabel metal2 s 326774 -960 326886 480 0 FreeSans 560 90 0 0 la_oenb[56]
port 479 nsew
flabel metal2 s 330362 -960 330474 480 0 FreeSans 560 90 0 0 la_oenb[57]
port 480 nsew
flabel metal2 s 333858 -960 333970 480 0 FreeSans 560 90 0 0 la_oenb[58]
port 481 nsew
flabel metal2 s 337446 -960 337558 480 0 FreeSans 560 90 0 0 la_oenb[59]
port 482 nsew
flabel metal2 s 145902 -960 146014 480 0 FreeSans 560 90 0 0 la_oenb[5]
port 483 nsew
flabel metal2 s 340942 -960 341054 480 0 FreeSans 560 90 0 0 la_oenb[60]
port 484 nsew
flabel metal2 s 344530 -960 344642 480 0 FreeSans 560 90 0 0 la_oenb[61]
port 485 nsew
flabel metal2 s 348026 -960 348138 480 0 FreeSans 560 90 0 0 la_oenb[62]
port 486 nsew
flabel metal2 s 351614 -960 351726 480 0 FreeSans 560 90 0 0 la_oenb[63]
port 487 nsew
flabel metal2 s 355202 -960 355314 480 0 FreeSans 560 90 0 0 la_oenb[64]
port 488 nsew
flabel metal2 s 358698 -960 358810 480 0 FreeSans 560 90 0 0 la_oenb[65]
port 489 nsew
flabel metal2 s 362286 -960 362398 480 0 FreeSans 560 90 0 0 la_oenb[66]
port 490 nsew
flabel metal2 s 365782 -960 365894 480 0 FreeSans 560 90 0 0 la_oenb[67]
port 491 nsew
flabel metal2 s 369370 -960 369482 480 0 FreeSans 560 90 0 0 la_oenb[68]
port 492 nsew
flabel metal2 s 372866 -960 372978 480 0 FreeSans 560 90 0 0 la_oenb[69]
port 493 nsew
flabel metal2 s 149490 -960 149602 480 0 FreeSans 560 90 0 0 la_oenb[6]
port 494 nsew
flabel metal2 s 376454 -960 376566 480 0 FreeSans 560 90 0 0 la_oenb[70]
port 495 nsew
flabel metal2 s 379950 -960 380062 480 0 FreeSans 560 90 0 0 la_oenb[71]
port 496 nsew
flabel metal2 s 383538 -960 383650 480 0 FreeSans 560 90 0 0 la_oenb[72]
port 497 nsew
flabel metal2 s 387126 -960 387238 480 0 FreeSans 560 90 0 0 la_oenb[73]
port 498 nsew
flabel metal2 s 390622 -960 390734 480 0 FreeSans 560 90 0 0 la_oenb[74]
port 499 nsew
flabel metal2 s 394210 -960 394322 480 0 FreeSans 560 90 0 0 la_oenb[75]
port 500 nsew
flabel metal2 s 397706 -960 397818 480 0 FreeSans 560 90 0 0 la_oenb[76]
port 501 nsew
flabel metal2 s 401294 -960 401406 480 0 FreeSans 560 90 0 0 la_oenb[77]
port 502 nsew
flabel metal2 s 404790 -960 404902 480 0 FreeSans 560 90 0 0 la_oenb[78]
port 503 nsew
flabel metal2 s 408378 -960 408490 480 0 FreeSans 560 90 0 0 la_oenb[79]
port 504 nsew
flabel metal2 s 152986 -960 153098 480 0 FreeSans 560 90 0 0 la_oenb[7]
port 505 nsew
flabel metal2 s 411874 -960 411986 480 0 FreeSans 560 90 0 0 la_oenb[80]
port 506 nsew
flabel metal2 s 415462 -960 415574 480 0 FreeSans 560 90 0 0 la_oenb[81]
port 507 nsew
flabel metal2 s 418958 -960 419070 480 0 FreeSans 560 90 0 0 la_oenb[82]
port 508 nsew
flabel metal2 s 422546 -960 422658 480 0 FreeSans 560 90 0 0 la_oenb[83]
port 509 nsew
flabel metal2 s 426134 -960 426246 480 0 FreeSans 560 90 0 0 la_oenb[84]
port 510 nsew
flabel metal2 s 429630 -960 429742 480 0 FreeSans 560 90 0 0 la_oenb[85]
port 511 nsew
flabel metal2 s 433218 -960 433330 480 0 FreeSans 560 90 0 0 la_oenb[86]
port 512 nsew
flabel metal2 s 436714 -960 436826 480 0 FreeSans 560 90 0 0 la_oenb[87]
port 513 nsew
flabel metal2 s 440302 -960 440414 480 0 FreeSans 560 90 0 0 la_oenb[88]
port 514 nsew
flabel metal2 s 443798 -960 443910 480 0 FreeSans 560 90 0 0 la_oenb[89]
port 515 nsew
flabel metal2 s 156574 -960 156686 480 0 FreeSans 560 90 0 0 la_oenb[8]
port 516 nsew
flabel metal2 s 447386 -960 447498 480 0 FreeSans 560 90 0 0 la_oenb[90]
port 517 nsew
flabel metal2 s 450882 -960 450994 480 0 FreeSans 560 90 0 0 la_oenb[91]
port 518 nsew
flabel metal2 s 454470 -960 454582 480 0 FreeSans 560 90 0 0 la_oenb[92]
port 519 nsew
flabel metal2 s 458058 -960 458170 480 0 FreeSans 560 90 0 0 la_oenb[93]
port 520 nsew
flabel metal2 s 461554 -960 461666 480 0 FreeSans 560 90 0 0 la_oenb[94]
port 521 nsew
flabel metal2 s 465142 -960 465254 480 0 FreeSans 560 90 0 0 la_oenb[95]
port 522 nsew
flabel metal2 s 468638 -960 468750 480 0 FreeSans 560 90 0 0 la_oenb[96]
port 523 nsew
flabel metal2 s 472226 -960 472338 480 0 FreeSans 560 90 0 0 la_oenb[97]
port 524 nsew
flabel metal2 s 475722 -960 475834 480 0 FreeSans 560 90 0 0 la_oenb[98]
port 525 nsew
flabel metal2 s 479310 -960 479422 480 0 FreeSans 560 90 0 0 la_oenb[99]
port 526 nsew
flabel metal2 s 160070 -960 160182 480 0 FreeSans 560 90 0 0 la_oenb[9]
port 527 nsew
flabel metal2 s 579774 -960 579886 480 0 FreeSans 560 90 0 0 user_clock2
port 528 nsew
flabel metal2 s 580970 -960 581082 480 0 FreeSans 560 90 0 0 user_irq[0]
port 529 nsew
flabel metal2 s 582166 -960 582278 480 0 FreeSans 560 90 0 0 user_irq[1]
port 530 nsew
flabel metal2 s 583362 -960 583474 480 0 FreeSans 560 90 0 0 user_irq[2]
port 531 nsew
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 181794 -7654 182414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 145794 -7654 146414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 109794 -7654 110414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal4 s 549234 -7654 549854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 513234 -7654 513854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 477234 354980 477854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 441234 -7654 441854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 405234 -7654 405854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 369234 354980 369854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 333234 -7654 333854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 297234 -7654 297854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 261234 354980 261854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 225234 -7654 225854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 189234 -7654 189854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 153234 -7654 153854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 117234 -7654 117854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 81234 -7654 81854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 45234 -7654 45854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal4 s 556674 -7654 557294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 520674 -7654 521294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 484674 -7654 485294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 448674 -7654 449294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 412674 -7654 413294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 376674 -7654 377294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 340674 -7654 341294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 304674 -7654 305294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 268674 -7654 269294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 232674 -7654 233294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 196674 -7654 197294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 160674 -7654 161294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 124674 -7654 125294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 88674 -7654 89294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 52674 -7654 53294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal4 s 564114 -7654 564734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 528114 -7654 528734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 492114 354980 492734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 456114 -7654 456734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 420114 -7654 420734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 384114 354980 384734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 348114 -7654 348734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 312114 -7654 312734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 276114 -7654 276734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 240114 -7654 240734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 204114 -7654 204734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 168114 -7654 168734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 132114 -7654 132734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 96114 -7654 96734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 60114 -7654 60734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 24114 -7654 24734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal4 s 560394 -7654 561014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 524394 -7654 525014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 488394 -7654 489014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 452394 -7654 453014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 416394 -7654 417014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 380394 -7654 381014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 344394 -7654 345014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 308394 354980 309014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 272394 -7654 273014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 236394 -7654 237014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 200394 354980 201014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 164394 -7654 165014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 128394 -7654 129014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 92394 354980 93014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 56394 -7654 57014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 531834 -7654 532454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 495834 -7654 496454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 459834 -7654 460454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 423834 -7654 424454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 387834 -7654 388454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 351834 -7654 352454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 315834 -7654 316454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 279834 -7654 280454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 243834 -7654 244454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 207834 -7654 208454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 171834 -7654 172454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 135834 -7654 136454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 99834 -7654 100454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 63834 -7654 64454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 27834 -7654 28454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 545514 -7654 546134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 509514 -7654 510134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 473514 -7654 474134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 437514 -7654 438134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 401514 -7654 402134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 365514 -7654 366134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 329514 -7654 330134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 293514 -7654 294134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 257514 -7654 258134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 221514 -7654 222134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 185514 354980 186134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 149514 -7654 150134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 113514 -7654 114134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 77514 354980 78134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 41514 -7654 42134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal4 s 552954 -7654 553574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 516954 -7654 517574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 480954 -7654 481574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 444954 -7654 445574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 408954 -7654 409574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 372954 -7654 373574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 336954 -7654 337574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 300954 -7654 301574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 264954 -7654 265574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 228954 -7654 229574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 192954 -7654 193574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 156954 -7654 157574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 120954 -7654 121574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 84954 -7654 85574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 48954 -7654 49574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal2 s 542 -960 654 480 0 FreeSans 560 90 0 0 wb_clk_i
port 540 nsew
flabel metal2 s 1646 -960 1758 480 0 FreeSans 560 90 0 0 wb_rst_i
port 541 nsew
flabel metal2 s 2842 -960 2954 480 0 FreeSans 560 90 0 0 wbs_ack_o
port 542 nsew
flabel metal2 s 7626 -960 7738 480 0 FreeSans 560 90 0 0 wbs_adr_i[0]
port 543 nsew
flabel metal2 s 47830 -960 47942 480 0 FreeSans 560 90 0 0 wbs_adr_i[10]
port 544 nsew
flabel metal2 s 51326 -960 51438 480 0 FreeSans 560 90 0 0 wbs_adr_i[11]
port 545 nsew
flabel metal2 s 54914 -960 55026 480 0 FreeSans 560 90 0 0 wbs_adr_i[12]
port 546 nsew
flabel metal2 s 58410 -960 58522 480 0 FreeSans 560 90 0 0 wbs_adr_i[13]
port 547 nsew
flabel metal2 s 61998 -960 62110 480 0 FreeSans 560 90 0 0 wbs_adr_i[14]
port 548 nsew
flabel metal2 s 65494 -960 65606 480 0 FreeSans 560 90 0 0 wbs_adr_i[15]
port 549 nsew
flabel metal2 s 69082 -960 69194 480 0 FreeSans 560 90 0 0 wbs_adr_i[16]
port 550 nsew
flabel metal2 s 72578 -960 72690 480 0 FreeSans 560 90 0 0 wbs_adr_i[17]
port 551 nsew
flabel metal2 s 76166 -960 76278 480 0 FreeSans 560 90 0 0 wbs_adr_i[18]
port 552 nsew
flabel metal2 s 79662 -960 79774 480 0 FreeSans 560 90 0 0 wbs_adr_i[19]
port 553 nsew
flabel metal2 s 12318 -960 12430 480 0 FreeSans 560 90 0 0 wbs_adr_i[1]
port 554 nsew
flabel metal2 s 83250 -960 83362 480 0 FreeSans 560 90 0 0 wbs_adr_i[20]
port 555 nsew
flabel metal2 s 86838 -960 86950 480 0 FreeSans 560 90 0 0 wbs_adr_i[21]
port 556 nsew
flabel metal2 s 90334 -960 90446 480 0 FreeSans 560 90 0 0 wbs_adr_i[22]
port 557 nsew
flabel metal2 s 93922 -960 94034 480 0 FreeSans 560 90 0 0 wbs_adr_i[23]
port 558 nsew
flabel metal2 s 97418 -960 97530 480 0 FreeSans 560 90 0 0 wbs_adr_i[24]
port 559 nsew
flabel metal2 s 101006 -960 101118 480 0 FreeSans 560 90 0 0 wbs_adr_i[25]
port 560 nsew
flabel metal2 s 104502 -960 104614 480 0 FreeSans 560 90 0 0 wbs_adr_i[26]
port 561 nsew
flabel metal2 s 108090 -960 108202 480 0 FreeSans 560 90 0 0 wbs_adr_i[27]
port 562 nsew
flabel metal2 s 111586 -960 111698 480 0 FreeSans 560 90 0 0 wbs_adr_i[28]
port 563 nsew
flabel metal2 s 115174 -960 115286 480 0 FreeSans 560 90 0 0 wbs_adr_i[29]
port 564 nsew
flabel metal2 s 17010 -960 17122 480 0 FreeSans 560 90 0 0 wbs_adr_i[2]
port 565 nsew
flabel metal2 s 118762 -960 118874 480 0 FreeSans 560 90 0 0 wbs_adr_i[30]
port 566 nsew
flabel metal2 s 122258 -960 122370 480 0 FreeSans 560 90 0 0 wbs_adr_i[31]
port 567 nsew
flabel metal2 s 21794 -960 21906 480 0 FreeSans 560 90 0 0 wbs_adr_i[3]
port 568 nsew
flabel metal2 s 26486 -960 26598 480 0 FreeSans 560 90 0 0 wbs_adr_i[4]
port 569 nsew
flabel metal2 s 30074 -960 30186 480 0 FreeSans 560 90 0 0 wbs_adr_i[5]
port 570 nsew
flabel metal2 s 33570 -960 33682 480 0 FreeSans 560 90 0 0 wbs_adr_i[6]
port 571 nsew
flabel metal2 s 37158 -960 37270 480 0 FreeSans 560 90 0 0 wbs_adr_i[7]
port 572 nsew
flabel metal2 s 40654 -960 40766 480 0 FreeSans 560 90 0 0 wbs_adr_i[8]
port 573 nsew
flabel metal2 s 44242 -960 44354 480 0 FreeSans 560 90 0 0 wbs_adr_i[9]
port 574 nsew
flabel metal2 s 4038 -960 4150 480 0 FreeSans 560 90 0 0 wbs_cyc_i
port 575 nsew
flabel metal2 s 8730 -960 8842 480 0 FreeSans 560 90 0 0 wbs_dat_i[0]
port 576 nsew
flabel metal2 s 48934 -960 49046 480 0 FreeSans 560 90 0 0 wbs_dat_i[10]
port 577 nsew
flabel metal2 s 52522 -960 52634 480 0 FreeSans 560 90 0 0 wbs_dat_i[11]
port 578 nsew
flabel metal2 s 56018 -960 56130 480 0 FreeSans 560 90 0 0 wbs_dat_i[12]
port 579 nsew
flabel metal2 s 59606 -960 59718 480 0 FreeSans 560 90 0 0 wbs_dat_i[13]
port 580 nsew
flabel metal2 s 63194 -960 63306 480 0 FreeSans 560 90 0 0 wbs_dat_i[14]
port 581 nsew
flabel metal2 s 66690 -960 66802 480 0 FreeSans 560 90 0 0 wbs_dat_i[15]
port 582 nsew
flabel metal2 s 70278 -960 70390 480 0 FreeSans 560 90 0 0 wbs_dat_i[16]
port 583 nsew
flabel metal2 s 73774 -960 73886 480 0 FreeSans 560 90 0 0 wbs_dat_i[17]
port 584 nsew
flabel metal2 s 77362 -960 77474 480 0 FreeSans 560 90 0 0 wbs_dat_i[18]
port 585 nsew
flabel metal2 s 80858 -960 80970 480 0 FreeSans 560 90 0 0 wbs_dat_i[19]
port 586 nsew
flabel metal2 s 13514 -960 13626 480 0 FreeSans 560 90 0 0 wbs_dat_i[1]
port 587 nsew
flabel metal2 s 84446 -960 84558 480 0 FreeSans 560 90 0 0 wbs_dat_i[20]
port 588 nsew
flabel metal2 s 87942 -960 88054 480 0 FreeSans 560 90 0 0 wbs_dat_i[21]
port 589 nsew
flabel metal2 s 91530 -960 91642 480 0 FreeSans 560 90 0 0 wbs_dat_i[22]
port 590 nsew
flabel metal2 s 95118 -960 95230 480 0 FreeSans 560 90 0 0 wbs_dat_i[23]
port 591 nsew
flabel metal2 s 98614 -960 98726 480 0 FreeSans 560 90 0 0 wbs_dat_i[24]
port 592 nsew
flabel metal2 s 102202 -960 102314 480 0 FreeSans 560 90 0 0 wbs_dat_i[25]
port 593 nsew
flabel metal2 s 105698 -960 105810 480 0 FreeSans 560 90 0 0 wbs_dat_i[26]
port 594 nsew
flabel metal2 s 109286 -960 109398 480 0 FreeSans 560 90 0 0 wbs_dat_i[27]
port 595 nsew
flabel metal2 s 112782 -960 112894 480 0 FreeSans 560 90 0 0 wbs_dat_i[28]
port 596 nsew
flabel metal2 s 116370 -960 116482 480 0 FreeSans 560 90 0 0 wbs_dat_i[29]
port 597 nsew
flabel metal2 s 18206 -960 18318 480 0 FreeSans 560 90 0 0 wbs_dat_i[2]
port 598 nsew
flabel metal2 s 119866 -960 119978 480 0 FreeSans 560 90 0 0 wbs_dat_i[30]
port 599 nsew
flabel metal2 s 123454 -960 123566 480 0 FreeSans 560 90 0 0 wbs_dat_i[31]
port 600 nsew
flabel metal2 s 22990 -960 23102 480 0 FreeSans 560 90 0 0 wbs_dat_i[3]
port 601 nsew
flabel metal2 s 27682 -960 27794 480 0 FreeSans 560 90 0 0 wbs_dat_i[4]
port 602 nsew
flabel metal2 s 31270 -960 31382 480 0 FreeSans 560 90 0 0 wbs_dat_i[5]
port 603 nsew
flabel metal2 s 34766 -960 34878 480 0 FreeSans 560 90 0 0 wbs_dat_i[6]
port 604 nsew
flabel metal2 s 38354 -960 38466 480 0 FreeSans 560 90 0 0 wbs_dat_i[7]
port 605 nsew
flabel metal2 s 41850 -960 41962 480 0 FreeSans 560 90 0 0 wbs_dat_i[8]
port 606 nsew
flabel metal2 s 45438 -960 45550 480 0 FreeSans 560 90 0 0 wbs_dat_i[9]
port 607 nsew
flabel metal2 s 9926 -960 10038 480 0 FreeSans 560 90 0 0 wbs_dat_o[0]
port 608 nsew
flabel metal2 s 50130 -960 50242 480 0 FreeSans 560 90 0 0 wbs_dat_o[10]
port 609 nsew
flabel metal2 s 53718 -960 53830 480 0 FreeSans 560 90 0 0 wbs_dat_o[11]
port 610 nsew
flabel metal2 s 57214 -960 57326 480 0 FreeSans 560 90 0 0 wbs_dat_o[12]
port 611 nsew
flabel metal2 s 60802 -960 60914 480 0 FreeSans 560 90 0 0 wbs_dat_o[13]
port 612 nsew
flabel metal2 s 64298 -960 64410 480 0 FreeSans 560 90 0 0 wbs_dat_o[14]
port 613 nsew
flabel metal2 s 67886 -960 67998 480 0 FreeSans 560 90 0 0 wbs_dat_o[15]
port 614 nsew
flabel metal2 s 71474 -960 71586 480 0 FreeSans 560 90 0 0 wbs_dat_o[16]
port 615 nsew
flabel metal2 s 74970 -960 75082 480 0 FreeSans 560 90 0 0 wbs_dat_o[17]
port 616 nsew
flabel metal2 s 78558 -960 78670 480 0 FreeSans 560 90 0 0 wbs_dat_o[18]
port 617 nsew
flabel metal2 s 82054 -960 82166 480 0 FreeSans 560 90 0 0 wbs_dat_o[19]
port 618 nsew
flabel metal2 s 14710 -960 14822 480 0 FreeSans 560 90 0 0 wbs_dat_o[1]
port 619 nsew
flabel metal2 s 85642 -960 85754 480 0 FreeSans 560 90 0 0 wbs_dat_o[20]
port 620 nsew
flabel metal2 s 89138 -960 89250 480 0 FreeSans 560 90 0 0 wbs_dat_o[21]
port 621 nsew
flabel metal2 s 92726 -960 92838 480 0 FreeSans 560 90 0 0 wbs_dat_o[22]
port 622 nsew
flabel metal2 s 96222 -960 96334 480 0 FreeSans 560 90 0 0 wbs_dat_o[23]
port 623 nsew
flabel metal2 s 99810 -960 99922 480 0 FreeSans 560 90 0 0 wbs_dat_o[24]
port 624 nsew
flabel metal2 s 103306 -960 103418 480 0 FreeSans 560 90 0 0 wbs_dat_o[25]
port 625 nsew
flabel metal2 s 106894 -960 107006 480 0 FreeSans 560 90 0 0 wbs_dat_o[26]
port 626 nsew
flabel metal2 s 110482 -960 110594 480 0 FreeSans 560 90 0 0 wbs_dat_o[27]
port 627 nsew
flabel metal2 s 113978 -960 114090 480 0 FreeSans 560 90 0 0 wbs_dat_o[28]
port 628 nsew
flabel metal2 s 117566 -960 117678 480 0 FreeSans 560 90 0 0 wbs_dat_o[29]
port 629 nsew
flabel metal2 s 19402 -960 19514 480 0 FreeSans 560 90 0 0 wbs_dat_o[2]
port 630 nsew
flabel metal2 s 121062 -960 121174 480 0 FreeSans 560 90 0 0 wbs_dat_o[30]
port 631 nsew
flabel metal2 s 124650 -960 124762 480 0 FreeSans 560 90 0 0 wbs_dat_o[31]
port 632 nsew
flabel metal2 s 24186 -960 24298 480 0 FreeSans 560 90 0 0 wbs_dat_o[3]
port 633 nsew
flabel metal2 s 28878 -960 28990 480 0 FreeSans 560 90 0 0 wbs_dat_o[4]
port 634 nsew
flabel metal2 s 32374 -960 32486 480 0 FreeSans 560 90 0 0 wbs_dat_o[5]
port 635 nsew
flabel metal2 s 35962 -960 36074 480 0 FreeSans 560 90 0 0 wbs_dat_o[6]
port 636 nsew
flabel metal2 s 39550 -960 39662 480 0 FreeSans 560 90 0 0 wbs_dat_o[7]
port 637 nsew
flabel metal2 s 43046 -960 43158 480 0 FreeSans 560 90 0 0 wbs_dat_o[8]
port 638 nsew
flabel metal2 s 46634 -960 46746 480 0 FreeSans 560 90 0 0 wbs_dat_o[9]
port 639 nsew
flabel metal2 s 11122 -960 11234 480 0 FreeSans 560 90 0 0 wbs_sel_i[0]
port 640 nsew
flabel metal2 s 15906 -960 16018 480 0 FreeSans 560 90 0 0 wbs_sel_i[1]
port 641 nsew
flabel metal2 s 20598 -960 20710 480 0 FreeSans 560 90 0 0 wbs_sel_i[2]
port 642 nsew
flabel metal2 s 25290 -960 25402 480 0 FreeSans 560 90 0 0 wbs_sel_i[3]
port 643 nsew
flabel metal2 s 5234 -960 5346 480 0 FreeSans 560 90 0 0 wbs_stb_i
port 644 nsew
flabel metal2 s 6430 -960 6542 480 0 FreeSans 560 90 0 0 wbs_we_i
port 645 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
